
module command4Cycle ( ri, ao, _reset, ai, ro, l0, l1, l2 );
input  ri, ao, _reset;
output ai, ro, l0, l1, l2;
    wire n6, csc0, csc1, _X11, _X13, _X14, _X16, _X17, _X18, _X19, _X20, _X21, 
        _X22, _X23, n1, n2, n3, n4;
    and2_1 _U29 ( .x(_X21), .a(ri), .b(csc0) );
    and2_1 _U28 ( .x(_X20), .a(_X18), .b(_X19) );
    and2_1 _U18 ( .x(_X14), .a(l1), .b(csc1) );
    and2_1 _U17 ( .x(_X13), .a(l1), .b(_X19) );
    and2_1 _U32 ( .x(_X23), .a(ri), .b(csc1) );
    and2_1 _U23 ( .x(_X17), .a(n6), .b(csc0) );
    and2_1 _U22 ( .x(_X16), .a(n6), .b(_X19) );
    or3_2 _U33 ( .x(csc1), .a(_X22), .b(l0), .c(_X23) );
    and2_1 _U13 ( .x(_X11), .a(_X19), .b(l0) );
    or3i_1 U1 ( .x(n6), .a(n1), .b(_X17), .c(_X16) );
    or3i_1 U2 ( .x(csc0), .a(_X22), .b(_X21), .c(_X20) );
    inv_0 U4 ( .x(_X19), .a(ri) );
    nor2_0 U6 ( .x(ro), .a(_X19), .b(n2) );
    aoi21_1 U7 ( .x(n2), .a(_X18), .b(csc0), .c(ao) );
    aoi31_1 U8 ( .x(n3), .a(csc0), .b(n4), .c(csc1), .d(ao) );
    aoi22_1 U10 ( .x(ai), .a(n3), .b(n6), .c(csc0), .d(_X18) );
    inv_0 U12 ( .x(_X22), .a(l1) );
    inv_0 U13 ( .x(n4), .a(l0) );
    nor2i_1 U14 ( .x(n1), .a(_reset), .b(ao) );
    or3i_2 U15 ( .x(l1), .a(n1), .b(_X14), .c(_X13) );
    inv_1 U16 ( .x(l2), .a(_X18) );
    inv_2 U17 ( .x(_X18), .a(n6) );
    nand2i_2 U18 ( .x(l0), .a(_X11), .b(n1) );
endmodule


module matched_delay_tic_com ( x, a );
input  a;
output x;
    assign x = a;
endmodule


module response4Cycle ( ri, ao, _reset, ai, ro, l0, l1, l2, l3 );
input  ri, ao, _reset;
output ai, ro, l0, l1, l2, l3;
    wire n2, n3, n4, csc0, csc1, _X7, _X9, _X8, _X10, _reset__not, _X13, 
        csc2__reset, _X11, _X14, csc2, _X16, _X18, _X20, csc0__reset, _X21, 
        l3_csc0_reset, _X25, _X26, _X30, _X31, csc1__reset, _X36, _X35, _X37, 
        n5, n6, n7, n8, n9, n10;
    or2_2 _U44 ( .x(l3_csc0_reset), .a(_reset__not), .b(l3) );
    and2_1 _U22_4 ( .x(n4), .a(n3), .b(_X13) );
    and2_1 _U22_3 ( .x(n3), .a(n2), .b(csc0) );
    and2_1 _U24 ( .x(csc2__reset), .a(_reset), .b(csc2) );
    and2_1 _U41 ( .x(_X26), .a(csc0), .b(_X25) );
    and2_1 _U57 ( .x(csc1__reset), .a(_reset), .b(csc1) );
    and2_1 _U53 ( .x(_X35), .a(_X7), .b(csc2) );
    and2_1 _U54 ( .x(_X37), .a(_X36), .b(csc2) );
    and2_1 _U47 ( .x(_X31), .a(csc1), .b(_X30) );
    and3_1 _U16 ( .x(_X10), .a(ri), .b(_X9), .c(csc1) );
    and2_1 _U15 ( .x(_X8), .a(_X7), .b(l0) );
    and2_1 _U22_5 ( .x(_X14), .a(n4), .b(csc1) );
    and2_1 _U21 ( .x(_X11), .a(l1), .b(csc2__reset) );
    and2_1 _U28 ( .x(_X18), .a(l2), .b(_X16) );
    and2_1 _U33 ( .x(_X20), .a(_X7), .b(l3) );
    and2_1 _U34 ( .x(_X21), .a(csc0__reset), .b(l3) );
    oai222_1 U1 ( .x(ro), .a(_X13), .b(n5), .c(_reset__not), .d(n6), .e(csc1), 
        .f(csc0) );
    inv_0 U2 ( .x(_reset__not), .a(_reset) );
    oai21_1 U3 ( .x(csc2), .a(csc1__reset), .b(_X7), .c(n7) );
    nor2_0 U4 ( .x(_X36), .a(_X14), .b(_X11) );
    ao21_1 U7 ( .x(csc0), .a(n10), .b(n8), .c(_X26) );
    inv_0 U9 ( .x(_X25), .a(l3_csc0_reset) );
    and3i_1 U11 ( .x(n2), .a(ao), .b(ri), .c(csc2__reset) );
    oa21_1 U12 ( .x(ai), .a(l3), .b(_X9), .c(ro) );
    nor3_0 U13 ( .x(n6), .a(l3), .b(l1), .c(l2) );
    nand2_0 U15 ( .x(n5), .a(csc0), .b(_reset) );
    nor2_0 U16 ( .x(n7), .a(_X35), .b(_X37) );
    inv_0 U17 ( .x(n8), .a(ao) );
    inv_0 U18 ( .x(csc0__reset), .a(n5) );
    inv_0 U20 ( .x(_X9), .a(csc0) );
    inv_0 U22 ( .x(_X16), .a(csc2) );
    inv_0 U23 ( .x(_X30), .a(l2) );
    nand3i_0 U24 ( .x(n9), .a(csc1), .b(_X30), .c(_X7) );
    nand2i_2 U25 ( .x(csc1), .a(_X31), .b(ri) );
    nor2_1 U26 ( .x(_X7), .a(ao), .b(_reset__not) );
    ao21_2 U27 ( .x(l2), .a(_X16), .b(n8), .c(_X18) );
    inv_2 U28 ( .x(l1), .a(_X36) );
    or3i_2 U29 ( .x(l3), .a(n9), .b(_X20), .c(_X21) );
    inv_0 U30 ( .x(n10), .a(_X13) );
    inv_1 U31 ( .x(l0), .a(_X13) );
    nor2_1 U32 ( .x(_X13), .a(_X10), .b(_X8) );
endmodule


module matched_delay_tic_resp ( x, a );
input  a;
output x;
    assign x = a;
endmodule


module tic ( c_req, c_ack, c_we, c_addr, r_req, r_ack, data_in, data_out, 
    reset_b, mc_req, mc_we, mc_adr, mc_dat, mc_ack, mr_req, mr_dat, mr_ack );
input  [10:0] c_addr;
input  [7:0] data_in;
output [7:0] data_out;
output [31:0] mc_adr;
output [31:0] mc_dat;
input  [31:0] mr_dat;
input  c_req, c_we, r_ack, reset_b, mc_ack, mr_req;
output c_ack, r_req, mc_req, mc_we, mr_ack;
    wire \c_addr[10] , \c_addr[9] , \c_addr[8] , \c_addr[7] , \c_addr[6] , 
        \c_addr[5] , \c_addr[4] , \c_addr[3] , \c_addr[2] , \c_addr[1] , 
        \c_addr[0] , \data_in[7] , \data_in[6] , \data_in[5] , \data_in[4] , 
        \data_in[3] , \data_in[2] , \data_in[1] , \data_in[0] , wl0, wl1, wl2, 
        \s[3] , \s[2] , \s[1] , \s[0] , cwr, crr, wr_ack, w_r, _66_net_, rwr, 
        rrr, rd_ack, r_r, _67_net_, \covResp/nl , \covResp/ni , \covResp/nh , 
        \convCom/nl , \convCom/nh ;
    assign mc_we = c_we;
    assign \c_addr[10]  = c_addr[10];
    assign \c_addr[9]  = c_addr[9];
    assign \c_addr[8]  = c_addr[8];
    assign \c_addr[7]  = c_addr[7];
    assign \c_addr[6]  = c_addr[6];
    assign \c_addr[5]  = c_addr[5];
    assign \c_addr[4]  = c_addr[4];
    assign \c_addr[3]  = c_addr[3];
    assign \c_addr[2]  = c_addr[2];
    assign \c_addr[1]  = c_addr[1];
    assign \c_addr[0]  = c_addr[0];
    assign \data_in[7]  = data_in[7];
    assign \data_in[6]  = data_in[6];
    assign \data_in[5]  = data_in[5];
    assign \data_in[4]  = data_in[4];
    assign \data_in[3]  = data_in[3];
    assign \data_in[2]  = data_in[2];
    assign \data_in[1]  = data_in[1];
    assign \data_in[0]  = data_in[0];
    assign mc_adr[31] = \c_addr[10] ;
    assign mc_adr[30] = \c_addr[10] ;
    assign mc_adr[29] = 1'b0;
    assign mc_adr[28] = 1'b0;
    assign mc_adr[27] = 1'b0;
    assign mc_adr[26] = 1'b0;
    assign mc_adr[25] = 1'b0;
    assign mc_adr[24] = 1'b0;
    assign mc_adr[23] = 1'b0;
    assign mc_adr[22] = 1'b0;
    assign mc_adr[21] = 1'b0;
    assign mc_adr[20] = 1'b0;
    assign mc_adr[19] = 1'b0;
    assign mc_adr[18] = 1'b0;
    assign mc_adr[17] = 1'b0;
    assign mc_adr[16] = 1'b0;
    assign mc_adr[15] = 1'b0;
    assign mc_adr[14] = 1'b0;
    assign mc_adr[13] = 1'b0;
    assign mc_adr[12] = 1'b0;
    assign mc_adr[11] = \c_addr[9] ;
    assign mc_adr[10] = \c_addr[8] ;
    assign mc_adr[9] = \c_addr[7] ;
    assign mc_adr[8] = \c_addr[6] ;
    assign mc_adr[7] = \c_addr[5] ;
    assign mc_adr[6] = \c_addr[4] ;
    assign mc_adr[5] = \c_addr[3] ;
    assign mc_adr[4] = \c_addr[2] ;
    assign mc_adr[3] = \c_addr[1] ;
    assign mc_adr[2] = \c_addr[0] ;
    assign mc_adr[1] = 1'b0;
    assign mc_adr[0] = 1'b0;
    assign mc_dat[31] = \data_in[7] ;
    assign mc_dat[30] = \data_in[6] ;
    assign mc_dat[29] = \data_in[5] ;
    assign mc_dat[28] = \data_in[4] ;
    assign mc_dat[27] = \data_in[3] ;
    assign mc_dat[26] = \data_in[2] ;
    assign mc_dat[25] = \data_in[1] ;
    assign mc_dat[24] = \data_in[0] ;
    command4Cycle cc ( .ri(cwr), .ao(mc_ack), ._reset(reset_b), .ai(wr_ack), 
        .ro(w_r), .l0(wl0), .l1(wl1), .l2(wl2) );
    matched_delay_tic_com delCom ( .x(mc_req), .a(_66_net_) );
    response4Cycle rc ( .ri(rrr), .ao(r_ack), ._reset(reset_b), .ai(rd_ack), 
        .ro(r_r), .l0(\s[0] ), .l1(\s[1] ), .l2(\s[2] ), .l3(\s[3] ) );
    matched_delay_tic_resp delResp ( .x(r_req), .a(_67_net_) );
    inv_1 \covResp/Uih  ( .x(\covResp/nh ), .a(rwr) );
    inv_1 \covResp/Uil  ( .x(\covResp/nl ), .a(rrr) );
    inv_1 \convCom/Uih  ( .x(\convCom/nh ), .a(cwr) );
    inv_1 \convCom/Uil  ( .x(\convCom/nl ), .a(crr) );
    ao23_2 \covResp/Ucl/U1/U1  ( .x(rrr), .a(mr_req), .b(rrr), .c(mr_req), .d(
        \covResp/ni ), .e(\covResp/nh ) );
    ao23_2 \convCom/Ucl/U1/U1  ( .x(crr), .a(c_req), .b(crr), .c(c_req), .d(
        \covResp/ni ), .e(\convCom/nh ) );
    ao23_2 \convCom/Uch/U1/U1  ( .x(cwr), .a(c_req), .b(cwr), .c(c_req), .d(
        mc_we), .e(\convCom/nl ) );
    ao23_2 \covResp/Uch/U1/U1  ( .x(rwr), .a(mr_req), .b(rwr), .c(mr_req), .d(
        mc_we), .e(\covResp/nl ) );
    latn_2 \wd1_reg[7]  ( .q(mc_dat[15]), .d(\data_in[7] ), .g(wl1) );
    latn_2 \wd1_reg[6]  ( .q(mc_dat[14]), .d(\data_in[6] ), .g(wl1) );
    latn_2 \wd1_reg[5]  ( .q(mc_dat[13]), .d(\data_in[5] ), .g(wl1) );
    latn_2 \wd1_reg[4]  ( .q(mc_dat[12]), .d(\data_in[4] ), .g(wl1) );
    latn_2 \wd1_reg[3]  ( .q(mc_dat[11]), .d(\data_in[3] ), .g(wl1) );
    latn_2 \wd1_reg[2]  ( .q(mc_dat[10]), .d(\data_in[2] ), .g(wl1) );
    latn_2 \wd1_reg[1]  ( .q(mc_dat[9]), .d(\data_in[1] ), .g(wl1) );
    latn_2 \wd1_reg[0]  ( .q(mc_dat[8]), .d(\data_in[0] ), .g(wl1) );
    latn_1 \wd0_reg[6]  ( .q(mc_dat[6]), .d(\data_in[6] ), .g(wl0) );
    latn_1 \wd0_reg[7]  ( .q(mc_dat[7]), .d(\data_in[7] ), .g(wl0) );
    latn_1 \wd0_reg[2]  ( .q(mc_dat[2]), .d(\data_in[2] ), .g(wl0) );
    latn_1 \wd0_reg[5]  ( .q(mc_dat[5]), .d(\data_in[5] ), .g(wl0) );
    latn_1 \wd0_reg[1]  ( .q(mc_dat[1]), .d(\data_in[1] ), .g(wl0) );
    latn_2 \wd0_reg[4]  ( .q(mc_dat[4]), .d(\data_in[4] ), .g(wl0) );
    latn_2 \wd0_reg[3]  ( .q(mc_dat[3]), .d(\data_in[3] ), .g(wl0) );
    latn_2 \wd0_reg[0]  ( .q(mc_dat[0]), .d(\data_in[0] ), .g(wl0) );
    inv_0 U2 ( .x(\covResp/ni ), .a(mc_we) );
    or2_1 U3 ( .x(_67_net_), .a(r_r), .b(rwr) );
    ao21_1 U4 ( .x(mr_ack), .a(rwr), .b(r_ack), .c(rd_ack) );
    or2_1 U5 ( .x(_66_net_), .a(crr), .b(w_r) );
    ao21_1 U6 ( .x(c_ack), .a(crr), .b(mc_ack), .c(wr_ack) );
    mx4_1 U7 ( .x(data_out[0]), .d0(mr_dat[0]), .sl0(\s[0] ), .d1(mr_dat[8]), 
        .sl1(\s[1] ), .d2(mr_dat[16]), .sl2(\s[2] ), .d3(mr_dat[24]), .sl3(
        \s[3] ) );
    mx4_1 U8 ( .x(data_out[1]), .d0(mr_dat[1]), .sl0(\s[0] ), .d1(mr_dat[9]), 
        .sl1(\s[1] ), .d2(mr_dat[17]), .sl2(\s[2] ), .d3(mr_dat[25]), .sl3(
        \s[3] ) );
    mx4_1 U9 ( .x(data_out[2]), .d0(mr_dat[2]), .sl0(\s[0] ), .d1(mr_dat[10]), 
        .sl1(\s[1] ), .d2(mr_dat[18]), .sl2(\s[2] ), .d3(mr_dat[26]), .sl3(
        \s[3] ) );
    mx4_1 U10 ( .x(data_out[3]), .d0(mr_dat[3]), .sl0(\s[0] ), .d1(mr_dat[11]), 
        .sl1(\s[1] ), .d2(mr_dat[19]), .sl2(\s[2] ), .d3(mr_dat[27]), .sl3(
        \s[3] ) );
    mx4_1 U11 ( .x(data_out[4]), .d0(mr_dat[4]), .sl0(\s[0] ), .d1(mr_dat[12]), 
        .sl1(\s[1] ), .d2(mr_dat[20]), .sl2(\s[2] ), .d3(mr_dat[28]), .sl3(
        \s[3] ) );
    mx4_1 U12 ( .x(data_out[5]), .d0(mr_dat[5]), .sl0(\s[0] ), .d1(mr_dat[13]), 
        .sl1(\s[1] ), .d2(mr_dat[21]), .sl2(\s[2] ), .d3(mr_dat[29]), .sl3(
        \s[3] ) );
    mx4_1 U13 ( .x(data_out[6]), .d0(mr_dat[6]), .sl0(\s[0] ), .d1(mr_dat[14]), 
        .sl1(\s[1] ), .d2(mr_dat[22]), .sl2(\s[2] ), .d3(mr_dat[30]), .sl3(
        \s[3] ) );
    mx4_1 U14 ( .x(data_out[7]), .d0(\s[0] ), .sl0(mr_dat[7]), .d1(\s[1] ), 
        .sl1(mr_dat[15]), .d2(\s[2] ), .sl2(mr_dat[23]), .d3(\s[3] ), .sl3(
        mr_dat[31]) );
    latn_1 \wd2_reg[6]  ( .q(mc_dat[22]), .d(\data_in[6] ), .g(wl2) );
    latn_1 \wd2_reg[7]  ( .q(mc_dat[23]), .d(\data_in[7] ), .g(wl2) );
    latn_1 \wd2_reg[0]  ( .q(mc_dat[16]), .d(\data_in[0] ), .g(wl2) );
    latn_1 \wd2_reg[1]  ( .q(mc_dat[17]), .d(\data_in[1] ), .g(wl2) );
    latn_1 \wd2_reg[3]  ( .q(mc_dat[19]), .d(\data_in[3] ), .g(wl2) );
    latn_1 \wd2_reg[2]  ( .q(mc_dat[18]), .d(\data_in[2] ), .g(wl2) );
    latn_1 \wd2_reg[5]  ( .q(mc_dat[21]), .d(\data_in[5] ), .g(wl2) );
    latn_1 \wd2_reg[4]  ( .q(mc_dat[20]), .d(\data_in[4] ), .g(wl2) );
endmodule


module chain_router0 ( eop_i, d0_i, d1_i, d2_i, d3_i, ack_i, eop_ox, d0_ox, 
    d1_ox, d2_ox, d3_ox, ack_ox, eop_oy, d0_oy, d1_oy, d2_oy, d3_oy, ack_oy, 
    nrst, test_si, test_se, test_so, phi1, phi2, phi3 );
input  eop_i, d0_i, d1_i, d2_i, d3_i, ack_ox, ack_oy, nrst, test_si, test_se, 
    phi1, phi2, phi3;
output ack_i, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, eop_oy, d0_oy, d1_oy, d2_oy, 
    d3_oy, test_so;
    wire \scan[2] , \scan[3] , ackx_l, nack_x, sx, acky_l, nack_y, sy, 
        \scan[0] , qa, qa_l, nroutex, routeAckx, nrouteAckx, qx, nqx, neopxy, 
        \scan[1] , sx_pl, nroutey, routeAcky, nrouteAcky, qy, nqy, sy_pl, rst, 
        n10, n11, n12, n1, n2, n3, n4, n5, n6, n7, n8, \cy/__tmp99/nr , 
        \cy/__tmp99/nd , \cx/__tmp99/nr , \cx/__tmp99/nd , \cye/nr , \cye/nd , 
        \cye/n2 , \cy3/__tmp99/loop , \cy2/__tmp99/loop , \cy1/__tmp99/loop , 
        \cy0/__tmp99/loop , \cxe/nr , \cxe/nd , \cxe/n2 , \cx3/__tmp99/loop , 
        \cx2/__tmp99/loop , \cx1/__tmp99/loop , \cx0/__tmp99/loop , 
        \sl_sy/l1_q , \sl_sy/mxl/muxout , \sl_sx/l1_q , \sl_sx/mxl/muxout , 
        \sl_qa/l1_q , \sl_qa/mxl/muxout , \slAcky/l1_q , \slAcky/mxl/muxout , 
        \slAckx/l1_q , \slAckx/mxl/muxout ;
    inv_1 U0 ( .x(rst), .a(nrst) );
    nor2_2 U5 ( .x(nack_x), .a(ackx_l), .b(rst) );
    nor2_2 U4 ( .x(nack_y), .a(acky_l), .b(rst) );
    nand4_1 U1 ( .x(ack_i), .a(n10), .b(n11), .c(n12), .d(neopxy) );
    and4_1 U8 ( .x(n10), .a(n1), .b(n2), .c(n3), .d(n4) );
    inv_1 U10 ( .x(n1), .a(d0_oy) );
    inv_1 U11 ( .x(n2), .a(d1_oy) );
    inv_1 U14 ( .x(n3), .a(d2_oy) );
    inv_1 U16 ( .x(n4), .a(d3_oy) );
    and4_1 U9 ( .x(n11), .a(n5), .b(n6), .c(n7), .d(n8) );
    inv_1 U17 ( .x(n5), .a(d0_ox) );
    inv_1 U18 ( .x(n6), .a(d1_ox) );
    inv_1 U19 ( .x(n7), .a(d2_ox) );
    inv_1 U20 ( .x(n8), .a(d3_ox) );
    nor2_1 U7 ( .x(n12), .a(nrouteAckx), .b(nrouteAcky) );
    nor2_1 U6 ( .x(neopxy), .a(eop_oy), .b(eop_ox) );
    nor2_1 U3 ( .x(nroutex), .a(d3_i), .b(d1_i) );
    nor2_1 U2 ( .x(nroutey), .a(d2_i), .b(d0_i) );
    nand2_1 U12 ( .x(qa), .a(nqx), .b(nqy) );
    nor2i_1 U15 ( .x(sx_pl), .a(qx), .b(nrouteAckx) );
    nor2i_1 U13 ( .x(sy_pl), .a(qy), .b(nrouteAcky) );
    inv_1 \cy/U1  ( .x(nrouteAcky), .a(routeAcky) );
    nor2_1 \cy/__tmp99/U1  ( .x(\cy/__tmp99/nr ), .a(nroutey), .b(qa_l) );
    nand2_1 \cy/__tmp99/U2  ( .x(\cy/__tmp99/nd ), .a(nroutey), .b(qa_l) );
    oai211_1 \cy/__tmp99/U3  ( .x(routeAcky), .a(nrouteAcky), .b(
        \cy/__tmp99/nr ), .c(\cy/__tmp99/nd ), .d(nrst) );
    inv_1 \cx/U1  ( .x(nrouteAckx), .a(routeAckx) );
    nor2_1 \cx/__tmp99/U1  ( .x(\cx/__tmp99/nr ), .a(nroutex), .b(qa_l) );
    nand2_1 \cx/__tmp99/U2  ( .x(\cx/__tmp99/nd ), .a(nroutex), .b(qa_l) );
    oai211_1 \cx/__tmp99/U3  ( .x(routeAckx), .a(nrouteAckx), .b(
        \cx/__tmp99/nr ), .c(\cx/__tmp99/nd ), .d(nrst) );
    nor3_1 \cye/Unr  ( .x(\cye/nr ), .a(eop_i), .b(nack_y), .c(sy) );
    nand3_1 \cye/Und  ( .x(\cye/nd ), .a(eop_i), .b(nack_y), .c(sy) );
    oa21_1 \cye/U1  ( .x(\cye/n2 ), .a(\cye/n2 ), .b(\cye/nr ), .c(\cye/nd )
         );
    inv_1 \cye/U3  ( .x(eop_oy), .a(\cye/n2 ) );
    ao31_1 \cy3/__tmp99/aoi  ( .x(\cy3/__tmp99/loop ), .a(d3_i), .b(nack_y), 
        .c(sy), .d(d3_oy) );
    ao31_1 \cy2/__tmp99/aoi  ( .x(\cy2/__tmp99/loop ), .a(d2_i), .b(nack_y), 
        .c(sy), .d(d2_oy) );
    ao31_1 \cy1/__tmp99/aoi  ( .x(\cy1/__tmp99/loop ), .a(d1_i), .b(nack_y), 
        .c(sy), .d(d1_oy) );
    ao31_1 \cy0/__tmp99/aoi  ( .x(\cy0/__tmp99/loop ), .a(d0_i), .b(nack_y), 
        .c(sy), .d(d0_oy) );
    nor3_1 \cxe/Unr  ( .x(\cxe/nr ), .a(eop_i), .b(nack_x), .c(sx) );
    nand3_1 \cxe/Und  ( .x(\cxe/nd ), .a(eop_i), .b(nack_x), .c(sx) );
    oa21_1 \cxe/U1  ( .x(\cxe/n2 ), .a(\cxe/n2 ), .b(\cxe/nr ), .c(\cxe/nd )
         );
    inv_1 \cxe/U3  ( .x(eop_ox), .a(\cxe/n2 ) );
    ao31_1 \cx3/__tmp99/aoi  ( .x(\cx3/__tmp99/loop ), .a(d3_i), .b(nack_x), 
        .c(sx), .d(d3_ox) );
    oa21_1 \cx3/__tmp99/outGate  ( .x(d3_ox), .a(d3_i), .b(nack_x), .c(
        \cx3/__tmp99/loop ) );
    ao31_1 \cx2/__tmp99/aoi  ( .x(\cx2/__tmp99/loop ), .a(d2_i), .b(nack_x), 
        .c(sx), .d(d2_ox) );
    oa21_1 \cx2/__tmp99/outGate  ( .x(d2_ox), .a(d2_i), .b(nack_x), .c(
        \cx2/__tmp99/loop ) );
    ao31_1 \cx1/__tmp99/aoi  ( .x(\cx1/__tmp99/loop ), .a(d1_i), .b(nack_x), 
        .c(sx), .d(d1_ox) );
    oa21_1 \cx1/__tmp99/outGate  ( .x(d1_ox), .a(d1_i), .b(nack_x), .c(
        \cx1/__tmp99/loop ) );
    ao31_1 \cx0/__tmp99/aoi  ( .x(\cx0/__tmp99/loop ), .a(d0_i), .b(nack_x), 
        .c(sx), .d(d0_ox) );
    oa21_1 \cx0/__tmp99/outGate  ( .x(d0_ox), .a(d0_i), .b(nack_x), .c(
        \cx0/__tmp99/loop ) );
    nand3_1 \sry/i0  ( .x(nqy), .a(neopxy), .b(nrst), .c(qy) );
    nand2_1 \sry/i1  ( .x(qy), .a(routeAcky), .b(nqy) );
    nand3_1 \srx/i0  ( .x(nqx), .a(neopxy), .b(nrst), .c(qx) );
    nand2_1 \srx/i1  ( .x(qx), .a(routeAckx), .b(nqx) );
    latn_1 \sl_sy/lph3  ( .q(sy), .d(\sl_sy/l1_q ), .g(phi3) );
    latn_1 \sl_sy/lph2  ( .q(\scan[2] ), .d(\sl_sy/l1_q ), .g(phi2) );
    mux2_1 \sl_sy/mxl/mux  ( .x(\sl_sy/mxl/muxout ), .d0(sy_pl), .sl(test_se), 
        .d1(\scan[1] ) );
    latn_1 \sl_sy/mxl/lph1  ( .q(\sl_sy/l1_q ), .d(\sl_sy/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_sx/lph3  ( .q(sx), .d(\sl_sx/l1_q ), .g(phi3) );
    latn_1 \sl_sx/lph2  ( .q(\scan[1] ), .d(\sl_sx/l1_q ), .g(phi2) );
    mux2_1 \sl_sx/mxl/mux  ( .x(\sl_sx/mxl/muxout ), .d0(sx_pl), .sl(test_se), 
        .d1(\scan[0] ) );
    latn_1 \sl_sx/mxl/lph1  ( .q(\sl_sx/l1_q ), .d(\sl_sx/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_qa/lph3  ( .q(qa_l), .d(\sl_qa/l1_q ), .g(phi3) );
    latn_1 \sl_qa/lph2  ( .q(\scan[0] ), .d(\sl_qa/l1_q ), .g(phi2) );
    mux2_1 \sl_qa/mxl/mux  ( .x(\sl_qa/mxl/muxout ), .d0(qa), .sl(test_se), 
        .d1(test_si) );
    latn_1 \sl_qa/mxl/lph1  ( .q(\sl_qa/l1_q ), .d(\sl_qa/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAcky/lph3  ( .q(acky_l), .d(\slAcky/l1_q ), .g(phi3) );
    latn_1 \slAcky/lph2  ( .q(test_so), .d(\slAcky/l1_q ), .g(phi2) );
    mux2_1 \slAcky/mxl/mux  ( .x(\slAcky/mxl/muxout ), .d0(ack_oy), .sl(
        test_se), .d1(\scan[3] ) );
    latn_1 \slAcky/mxl/lph1  ( .q(\slAcky/l1_q ), .d(\slAcky/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAckx/lph3  ( .q(ackx_l), .d(\slAckx/l1_q ), .g(phi3) );
    latn_1 \slAckx/lph2  ( .q(\scan[3] ), .d(\slAckx/l1_q ), .g(phi2) );
    mux2_1 \slAckx/mxl/mux  ( .x(\slAckx/mxl/muxout ), .d0(ack_ox), .sl(
        test_se), .d1(\scan[2] ) );
    latn_1 \slAckx/mxl/lph1  ( .q(\slAckx/l1_q ), .d(\slAckx/mxl/muxout ), .g(
        phi1) );
    oa21_2 U21 ( .x(d2_oy), .a(d2_i), .b(nack_y), .c(\cy2/__tmp99/loop ) );
    oa21_2 U22 ( .x(d1_oy), .a(d1_i), .b(nack_y), .c(\cy1/__tmp99/loop ) );
    oa21_2 U23 ( .x(d3_oy), .a(d3_i), .b(nack_y), .c(\cy3/__tmp99/loop ) );
    oa21_2 U24 ( .x(d0_oy), .a(d0_i), .b(nack_y), .c(\cy0/__tmp99/loop ) );
endmodule


module chain_router1 ( eop_i, d0_i, d1_i, d2_i, d3_i, ack_i, eop_ox, d0_ox, 
    d1_ox, d2_ox, d3_ox, ack_ox, eop_oy, d0_oy, d1_oy, d2_oy, d3_oy, ack_oy, 
    nrst, test_si, test_se, test_so, phi1, phi2, phi3 );
input  eop_i, d0_i, d1_i, d2_i, d3_i, ack_ox, ack_oy, nrst, test_si, test_se, 
    phi1, phi2, phi3;
output ack_i, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, eop_oy, d0_oy, d1_oy, d2_oy, 
    d3_oy, test_so;
    wire \scan[2] , \scan[3] , ackx_l, nack_x, sx, acky_l, nack_y, sy, 
        \scan[0] , qa, qa_l, nroutex, routeAckx, nrouteAckx, qx, nqx, neopxy, 
        \scan[1] , sx_pl, nroutey, routeAcky, nrouteAcky, qy, nqy, sy_pl, rst, 
        n10, n11, n12, n1, n2, n3, n4, n5, n6, n7, n8, \cy/__tmp99/nr , 
        \cy/__tmp99/nd , \cx/__tmp99/nr , \cx/__tmp99/nd , \cye/nr , \cye/nd , 
        \cye/n2 , \cy3/__tmp99/loop , \cy2/__tmp99/loop , \cy1/__tmp99/loop , 
        \cy0/__tmp99/loop , \cxe/nr , \cxe/nd , \cxe/n2 , \cx3/__tmp99/loop , 
        \cx2/__tmp99/loop , \cx1/__tmp99/loop , \cx0/__tmp99/loop , 
        \sl_sy/l1_q , \sl_sy/mxl/muxout , \sl_sx/l1_q , \sl_sx/mxl/muxout , 
        \sl_qa/l1_q , \sl_qa/mxl/muxout , \slAcky/l1_q , \slAcky/mxl/muxout , 
        \slAckx/l1_q , \slAckx/mxl/muxout ;
    inv_1 U0 ( .x(rst), .a(nrst) );
    nor2_2 U5 ( .x(nack_x), .a(ackx_l), .b(rst) );
    nor2_2 U4 ( .x(nack_y), .a(acky_l), .b(rst) );
    nand4_1 U1 ( .x(ack_i), .a(n10), .b(n11), .c(n12), .d(neopxy) );
    and4_1 U8 ( .x(n10), .a(n1), .b(n2), .c(n3), .d(n4) );
    inv_1 U10 ( .x(n1), .a(d0_oy) );
    inv_1 U11 ( .x(n2), .a(d1_oy) );
    inv_1 U14 ( .x(n3), .a(d2_oy) );
    inv_1 U16 ( .x(n4), .a(d3_oy) );
    and4_1 U9 ( .x(n11), .a(n5), .b(n6), .c(n7), .d(n8) );
    inv_1 U17 ( .x(n5), .a(d0_ox) );
    inv_1 U18 ( .x(n6), .a(d1_ox) );
    inv_1 U19 ( .x(n7), .a(d2_ox) );
    inv_1 U20 ( .x(n8), .a(d3_ox) );
    nor2_1 U7 ( .x(n12), .a(nrouteAckx), .b(nrouteAcky) );
    nor2_1 U6 ( .x(neopxy), .a(eop_oy), .b(eop_ox) );
    nor2_1 U3 ( .x(nroutex), .a(d3_i), .b(d1_i) );
    nor2_1 U2 ( .x(nroutey), .a(d2_i), .b(d0_i) );
    nand2_1 U12 ( .x(qa), .a(nqx), .b(nqy) );
    nor2i_1 U15 ( .x(sx_pl), .a(qx), .b(nrouteAckx) );
    nor2i_1 U13 ( .x(sy_pl), .a(qy), .b(nrouteAcky) );
    inv_1 \cy/U1  ( .x(nrouteAcky), .a(routeAcky) );
    nor2_1 \cy/__tmp99/U1  ( .x(\cy/__tmp99/nr ), .a(nroutey), .b(qa_l) );
    nand2_1 \cy/__tmp99/U2  ( .x(\cy/__tmp99/nd ), .a(nroutey), .b(qa_l) );
    oai211_1 \cy/__tmp99/U3  ( .x(routeAcky), .a(nrouteAcky), .b(
        \cy/__tmp99/nr ), .c(\cy/__tmp99/nd ), .d(nrst) );
    inv_1 \cx/U1  ( .x(nrouteAckx), .a(routeAckx) );
    nor2_1 \cx/__tmp99/U1  ( .x(\cx/__tmp99/nr ), .a(nroutex), .b(qa_l) );
    nand2_1 \cx/__tmp99/U2  ( .x(\cx/__tmp99/nd ), .a(nroutex), .b(qa_l) );
    oai211_1 \cx/__tmp99/U3  ( .x(routeAckx), .a(nrouteAckx), .b(
        \cx/__tmp99/nr ), .c(\cx/__tmp99/nd ), .d(nrst) );
    nor3_1 \cye/Unr  ( .x(\cye/nr ), .a(eop_i), .b(nack_y), .c(sy) );
    nand3_1 \cye/Und  ( .x(\cye/nd ), .a(eop_i), .b(nack_y), .c(sy) );
    oa21_1 \cye/U1  ( .x(\cye/n2 ), .a(\cye/n2 ), .b(\cye/nr ), .c(\cye/nd )
         );
    inv_1 \cye/U3  ( .x(eop_oy), .a(\cye/n2 ) );
    ao31_1 \cy3/__tmp99/aoi  ( .x(\cy3/__tmp99/loop ), .a(d3_i), .b(nack_y), 
        .c(sy), .d(d3_oy) );
    oa21_1 \cy3/__tmp99/outGate  ( .x(d3_oy), .a(d3_i), .b(nack_y), .c(
        \cy3/__tmp99/loop ) );
    ao31_1 \cy2/__tmp99/aoi  ( .x(\cy2/__tmp99/loop ), .a(d2_i), .b(nack_y), 
        .c(sy), .d(d2_oy) );
    oa21_1 \cy2/__tmp99/outGate  ( .x(d2_oy), .a(d2_i), .b(nack_y), .c(
        \cy2/__tmp99/loop ) );
    ao31_1 \cy1/__tmp99/aoi  ( .x(\cy1/__tmp99/loop ), .a(d1_i), .b(nack_y), 
        .c(sy), .d(d1_oy) );
    oa21_1 \cy1/__tmp99/outGate  ( .x(d1_oy), .a(d1_i), .b(nack_y), .c(
        \cy1/__tmp99/loop ) );
    ao31_1 \cy0/__tmp99/aoi  ( .x(\cy0/__tmp99/loop ), .a(d0_i), .b(nack_y), 
        .c(sy), .d(d0_oy) );
    oa21_1 \cy0/__tmp99/outGate  ( .x(d0_oy), .a(d0_i), .b(nack_y), .c(
        \cy0/__tmp99/loop ) );
    nor3_1 \cxe/Unr  ( .x(\cxe/nr ), .a(eop_i), .b(nack_x), .c(sx) );
    nand3_1 \cxe/Und  ( .x(\cxe/nd ), .a(eop_i), .b(nack_x), .c(sx) );
    oa21_1 \cxe/U1  ( .x(\cxe/n2 ), .a(\cxe/n2 ), .b(\cxe/nr ), .c(\cxe/nd )
         );
    inv_1 \cxe/U3  ( .x(eop_ox), .a(\cxe/n2 ) );
    ao31_1 \cx3/__tmp99/aoi  ( .x(\cx3/__tmp99/loop ), .a(d3_i), .b(nack_x), 
        .c(sx), .d(d3_ox) );
    oa21_1 \cx3/__tmp99/outGate  ( .x(d3_ox), .a(d3_i), .b(nack_x), .c(
        \cx3/__tmp99/loop ) );
    ao31_1 \cx2/__tmp99/aoi  ( .x(\cx2/__tmp99/loop ), .a(d2_i), .b(nack_x), 
        .c(sx), .d(d2_ox) );
    oa21_1 \cx2/__tmp99/outGate  ( .x(d2_ox), .a(d2_i), .b(nack_x), .c(
        \cx2/__tmp99/loop ) );
    ao31_1 \cx1/__tmp99/aoi  ( .x(\cx1/__tmp99/loop ), .a(d1_i), .b(nack_x), 
        .c(sx), .d(d1_ox) );
    oa21_1 \cx1/__tmp99/outGate  ( .x(d1_ox), .a(d1_i), .b(nack_x), .c(
        \cx1/__tmp99/loop ) );
    ao31_1 \cx0/__tmp99/aoi  ( .x(\cx0/__tmp99/loop ), .a(d0_i), .b(nack_x), 
        .c(sx), .d(d0_ox) );
    oa21_1 \cx0/__tmp99/outGate  ( .x(d0_ox), .a(d0_i), .b(nack_x), .c(
        \cx0/__tmp99/loop ) );
    nand3_1 \sry/i0  ( .x(nqy), .a(neopxy), .b(nrst), .c(qy) );
    nand2_1 \sry/i1  ( .x(qy), .a(routeAcky), .b(nqy) );
    nand3_1 \srx/i0  ( .x(nqx), .a(neopxy), .b(nrst), .c(qx) );
    nand2_1 \srx/i1  ( .x(qx), .a(routeAckx), .b(nqx) );
    latn_1 \sl_sy/lph3  ( .q(sy), .d(\sl_sy/l1_q ), .g(phi3) );
    latn_1 \sl_sy/lph2  ( .q(\scan[2] ), .d(\sl_sy/l1_q ), .g(phi2) );
    mux2_1 \sl_sy/mxl/mux  ( .x(\sl_sy/mxl/muxout ), .d0(sy_pl), .sl(test_se), 
        .d1(\scan[1] ) );
    latn_1 \sl_sy/mxl/lph1  ( .q(\sl_sy/l1_q ), .d(\sl_sy/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_sx/lph3  ( .q(sx), .d(\sl_sx/l1_q ), .g(phi3) );
    latn_1 \sl_sx/lph2  ( .q(\scan[1] ), .d(\sl_sx/l1_q ), .g(phi2) );
    mux2_1 \sl_sx/mxl/mux  ( .x(\sl_sx/mxl/muxout ), .d0(sx_pl), .sl(test_se), 
        .d1(\scan[0] ) );
    latn_1 \sl_sx/mxl/lph1  ( .q(\sl_sx/l1_q ), .d(\sl_sx/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_qa/lph3  ( .q(qa_l), .d(\sl_qa/l1_q ), .g(phi3) );
    latn_1 \sl_qa/lph2  ( .q(\scan[0] ), .d(\sl_qa/l1_q ), .g(phi2) );
    mux2_1 \sl_qa/mxl/mux  ( .x(\sl_qa/mxl/muxout ), .d0(qa), .sl(test_se), 
        .d1(test_si) );
    latn_1 \sl_qa/mxl/lph1  ( .q(\sl_qa/l1_q ), .d(\sl_qa/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAcky/lph3  ( .q(acky_l), .d(\slAcky/l1_q ), .g(phi3) );
    latn_1 \slAcky/lph2  ( .q(test_so), .d(\slAcky/l1_q ), .g(phi2) );
    mux2_1 \slAcky/mxl/mux  ( .x(\slAcky/mxl/muxout ), .d0(ack_oy), .sl(
        test_se), .d1(\scan[3] ) );
    latn_1 \slAcky/mxl/lph1  ( .q(\slAcky/l1_q ), .d(\slAcky/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAckx/lph3  ( .q(ackx_l), .d(\slAckx/l1_q ), .g(phi3) );
    latn_1 \slAckx/lph2  ( .q(\scan[3] ), .d(\slAckx/l1_q ), .g(phi2) );
    mux2_1 \slAckx/mxl/mux  ( .x(\slAckx/mxl/muxout ), .d0(ack_ox), .sl(
        test_se), .d1(\scan[2] ) );
    latn_1 \slAckx/mxl/lph1  ( .q(\slAckx/l1_q ), .d(\slAckx/mxl/muxout ), .g(
        phi1) );
endmodule


module chain_router2 ( eop_i, d0_i, d1_i, d2_i, d3_i, ack_i, eop_ox, d0_ox, 
    d1_ox, d2_ox, d3_ox, ack_ox, eop_oy, d0_oy, d1_oy, d2_oy, d3_oy, ack_oy, 
    nrst, test_si, test_se, test_so, phi1, phi2, phi3 );
input  eop_i, d0_i, d1_i, d2_i, d3_i, ack_ox, ack_oy, nrst, test_si, test_se, 
    phi1, phi2, phi3;
output ack_i, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, eop_oy, d0_oy, d1_oy, d2_oy, 
    d3_oy, test_so;
    wire \scan[2] , \scan[3] , ackx_l, nack_x, sx, acky_l, nack_y, sy, 
        \scan[0] , qa, qa_l, nroutex, routeAckx, nrouteAckx, qx, nqx, neopxy, 
        \scan[1] , sx_pl, nroutey, routeAcky, nrouteAcky, qy, nqy, sy_pl, rst, 
        n10, n11, n12, n1, n2, n3, n4, n5, n6, n7, n8, \cy/__tmp99/nr , 
        \cy/__tmp99/nd , \cx/__tmp99/nr , \cx/__tmp99/nd , \cye/nr , \cye/nd , 
        \cye/n2 , \cy3/__tmp99/loop , \cy2/__tmp99/loop , \cy1/__tmp99/loop , 
        \cy0/__tmp99/loop , \cxe/nr , \cxe/nd , \cxe/n2 , \cx3/__tmp99/loop , 
        \cx2/__tmp99/loop , \cx1/__tmp99/loop , \cx0/__tmp99/loop , 
        \sl_sy/l1_q , \sl_sy/mxl/muxout , \sl_sx/l1_q , \sl_sx/mxl/muxout , 
        \sl_qa/l1_q , \sl_qa/mxl/muxout , \slAcky/l1_q , \slAcky/mxl/muxout , 
        \slAckx/l1_q , \slAckx/mxl/muxout ;
    inv_1 U0 ( .x(rst), .a(nrst) );
    nor2_2 U5 ( .x(nack_x), .a(ackx_l), .b(rst) );
    nor2_2 U4 ( .x(nack_y), .a(acky_l), .b(rst) );
    nand4_1 U1 ( .x(ack_i), .a(n10), .b(n11), .c(n12), .d(neopxy) );
    and4_1 U8 ( .x(n10), .a(n1), .b(n2), .c(n3), .d(n4) );
    inv_1 U10 ( .x(n1), .a(d0_oy) );
    inv_1 U11 ( .x(n2), .a(d1_oy) );
    inv_1 U14 ( .x(n3), .a(d2_oy) );
    inv_1 U16 ( .x(n4), .a(d3_oy) );
    and4_1 U9 ( .x(n11), .a(n5), .b(n6), .c(n7), .d(n8) );
    inv_1 U17 ( .x(n5), .a(d0_ox) );
    inv_1 U18 ( .x(n6), .a(d1_ox) );
    inv_1 U19 ( .x(n7), .a(d2_ox) );
    inv_1 U20 ( .x(n8), .a(d3_ox) );
    nor2_1 U7 ( .x(n12), .a(nrouteAckx), .b(nrouteAcky) );
    nor2_1 U6 ( .x(neopxy), .a(eop_oy), .b(eop_ox) );
    nor2_1 U3 ( .x(nroutex), .a(d3_i), .b(d1_i) );
    nor2_1 U2 ( .x(nroutey), .a(d2_i), .b(d0_i) );
    nand2_1 U12 ( .x(qa), .a(nqx), .b(nqy) );
    nor2i_1 U15 ( .x(sx_pl), .a(qx), .b(nrouteAckx) );
    nor2i_1 U13 ( .x(sy_pl), .a(qy), .b(nrouteAcky) );
    inv_1 \cy/U1  ( .x(nrouteAcky), .a(routeAcky) );
    nor2_1 \cy/__tmp99/U1  ( .x(\cy/__tmp99/nr ), .a(nroutey), .b(qa_l) );
    nand2_1 \cy/__tmp99/U2  ( .x(\cy/__tmp99/nd ), .a(nroutey), .b(qa_l) );
    oai211_1 \cy/__tmp99/U3  ( .x(routeAcky), .a(nrouteAcky), .b(
        \cy/__tmp99/nr ), .c(\cy/__tmp99/nd ), .d(nrst) );
    inv_1 \cx/U1  ( .x(nrouteAckx), .a(routeAckx) );
    nor2_1 \cx/__tmp99/U1  ( .x(\cx/__tmp99/nr ), .a(nroutex), .b(qa_l) );
    nand2_1 \cx/__tmp99/U2  ( .x(\cx/__tmp99/nd ), .a(nroutex), .b(qa_l) );
    oai211_1 \cx/__tmp99/U3  ( .x(routeAckx), .a(nrouteAckx), .b(
        \cx/__tmp99/nr ), .c(\cx/__tmp99/nd ), .d(nrst) );
    nor3_1 \cye/Unr  ( .x(\cye/nr ), .a(eop_i), .b(nack_y), .c(sy) );
    nand3_1 \cye/Und  ( .x(\cye/nd ), .a(eop_i), .b(nack_y), .c(sy) );
    oa21_1 \cye/U1  ( .x(\cye/n2 ), .a(\cye/n2 ), .b(\cye/nr ), .c(\cye/nd )
         );
    inv_1 \cye/U3  ( .x(eop_oy), .a(\cye/n2 ) );
    ao31_1 \cy3/__tmp99/aoi  ( .x(\cy3/__tmp99/loop ), .a(d3_i), .b(nack_y), 
        .c(sy), .d(d3_oy) );
    ao31_1 \cy2/__tmp99/aoi  ( .x(\cy2/__tmp99/loop ), .a(d2_i), .b(nack_y), 
        .c(sy), .d(d2_oy) );
    ao31_1 \cy1/__tmp99/aoi  ( .x(\cy1/__tmp99/loop ), .a(d1_i), .b(nack_y), 
        .c(sy), .d(d1_oy) );
    ao31_1 \cy0/__tmp99/aoi  ( .x(\cy0/__tmp99/loop ), .a(d0_i), .b(nack_y), 
        .c(sy), .d(d0_oy) );
    nor3_1 \cxe/Unr  ( .x(\cxe/nr ), .a(eop_i), .b(nack_x), .c(sx) );
    nand3_1 \cxe/Und  ( .x(\cxe/nd ), .a(eop_i), .b(nack_x), .c(sx) );
    oa21_1 \cxe/U1  ( .x(\cxe/n2 ), .a(\cxe/n2 ), .b(\cxe/nr ), .c(\cxe/nd )
         );
    inv_1 \cxe/U3  ( .x(eop_ox), .a(\cxe/n2 ) );
    ao31_1 \cx3/__tmp99/aoi  ( .x(\cx3/__tmp99/loop ), .a(d3_i), .b(nack_x), 
        .c(sx), .d(d3_ox) );
    ao31_1 \cx2/__tmp99/aoi  ( .x(\cx2/__tmp99/loop ), .a(d2_i), .b(nack_x), 
        .c(sx), .d(d2_ox) );
    ao31_1 \cx1/__tmp99/aoi  ( .x(\cx1/__tmp99/loop ), .a(d1_i), .b(nack_x), 
        .c(sx), .d(d1_ox) );
    ao31_1 \cx0/__tmp99/aoi  ( .x(\cx0/__tmp99/loop ), .a(d0_i), .b(nack_x), 
        .c(sx), .d(d0_ox) );
    nand3_1 \sry/i0  ( .x(nqy), .a(neopxy), .b(nrst), .c(qy) );
    nand2_1 \sry/i1  ( .x(qy), .a(routeAcky), .b(nqy) );
    nand3_1 \srx/i0  ( .x(nqx), .a(neopxy), .b(nrst), .c(qx) );
    nand2_1 \srx/i1  ( .x(qx), .a(routeAckx), .b(nqx) );
    latn_1 \sl_sy/lph3  ( .q(sy), .d(\sl_sy/l1_q ), .g(phi3) );
    latn_1 \sl_sy/lph2  ( .q(\scan[2] ), .d(\sl_sy/l1_q ), .g(phi2) );
    mux2_1 \sl_sy/mxl/mux  ( .x(\sl_sy/mxl/muxout ), .d0(sy_pl), .sl(test_se), 
        .d1(\scan[1] ) );
    latn_1 \sl_sy/mxl/lph1  ( .q(\sl_sy/l1_q ), .d(\sl_sy/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_sx/lph3  ( .q(sx), .d(\sl_sx/l1_q ), .g(phi3) );
    latn_1 \sl_sx/lph2  ( .q(\scan[1] ), .d(\sl_sx/l1_q ), .g(phi2) );
    mux2_1 \sl_sx/mxl/mux  ( .x(\sl_sx/mxl/muxout ), .d0(sx_pl), .sl(test_se), 
        .d1(\scan[0] ) );
    latn_1 \sl_sx/mxl/lph1  ( .q(\sl_sx/l1_q ), .d(\sl_sx/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_qa/lph3  ( .q(qa_l), .d(\sl_qa/l1_q ), .g(phi3) );
    latn_1 \sl_qa/lph2  ( .q(\scan[0] ), .d(\sl_qa/l1_q ), .g(phi2) );
    mux2_1 \sl_qa/mxl/mux  ( .x(\sl_qa/mxl/muxout ), .d0(qa), .sl(test_se), 
        .d1(test_si) );
    latn_1 \sl_qa/mxl/lph1  ( .q(\sl_qa/l1_q ), .d(\sl_qa/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAcky/lph3  ( .q(acky_l), .d(\slAcky/l1_q ), .g(phi3) );
    latn_1 \slAcky/lph2  ( .q(test_so), .d(\slAcky/l1_q ), .g(phi2) );
    mux2_1 \slAcky/mxl/mux  ( .x(\slAcky/mxl/muxout ), .d0(ack_oy), .sl(
        test_se), .d1(\scan[3] ) );
    latn_1 \slAcky/mxl/lph1  ( .q(\slAcky/l1_q ), .d(\slAcky/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAckx/lph3  ( .q(ackx_l), .d(\slAckx/l1_q ), .g(phi3) );
    latn_1 \slAckx/lph2  ( .q(\scan[3] ), .d(\slAckx/l1_q ), .g(phi2) );
    mux2_1 \slAckx/mxl/mux  ( .x(\slAckx/mxl/muxout ), .d0(ack_ox), .sl(
        test_se), .d1(\scan[2] ) );
    latn_1 \slAckx/mxl/lph1  ( .q(\slAckx/l1_q ), .d(\slAckx/mxl/muxout ), .g(
        phi1) );
    oa21_2 U21 ( .x(d3_oy), .a(d3_i), .b(nack_y), .c(\cy3/__tmp99/loop ) );
    oa21_2 U22 ( .x(d2_oy), .a(d2_i), .b(nack_y), .c(\cy2/__tmp99/loop ) );
    oa21_2 U23 ( .x(d1_ox), .a(d1_i), .b(nack_x), .c(\cx1/__tmp99/loop ) );
    oa21_2 U24 ( .x(d3_ox), .a(d3_i), .b(nack_x), .c(\cx3/__tmp99/loop ) );
    oa21_2 U25 ( .x(d2_ox), .a(d2_i), .b(nack_x), .c(\cx2/__tmp99/loop ) );
    oa21_2 U26 ( .x(d0_oy), .a(d0_i), .b(nack_y), .c(\cy0/__tmp99/loop ) );
    oa21_2 U27 ( .x(d0_ox), .a(d0_i), .b(nack_x), .c(\cx0/__tmp99/loop ) );
    oa21_2 U28 ( .x(d1_oy), .a(d1_i), .b(nack_y), .c(\cy1/__tmp99/loop ) );
endmodule


module chain_arbiter0 ( eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, ack_ix, eop_iy, 
    d0_iy, d1_iy, d2_iy, d3_iy, ack_iy, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, 
    eop_oy, d0_oy, d1_oy, d2_oy, d3_oy, ack_oxy, rst, test_si, test_se, 
    test_so, phi1, phi2, phi3 );
input  eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, eop_iy, d0_iy, d1_iy, d2_iy, d3_iy, 
    ack_oxy, rst, test_si, test_se, phi1, phi2, phi3;
output ack_ix, ack_iy, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, eop_oy, d0_oy, 
    d1_oy, d2_oy, d3_oy, test_so;
    wire \scan[1] , \scan[2] , ackx_l, nack_x, sx, acky_l, nack_y, sy, mrx, 
        req_x, mry, req_y, gx, gy, \scan[0] , sx_pl, sy_pl, n1x, n2x, n1y, n2y, 
        n5x, n6x, n5y, n6y, \cye/nr , \cye/nd , \cye/n2 , \cy3/__tmp99/loop , 
        \cy2/__tmp99/loop , \cy1/__tmp99/loop , \cy0/__tmp99/loop , \cxe/nr , 
        \cxe/nd , \cxe/n2 , \cx3/__tmp99/loop , \cx2/__tmp99/loop , 
        \cx1/__tmp99/loop , \cx0/__tmp99/loop , \mtx/gr2 , \mtx/gr1 , \sry/qz , 
        \srx/qz , \sl_sy/l1_q , \sl_sy/mxl/muxout , \sl_sx/l1_q , 
        \sl_sx/mxl/muxout , \slAcky/l1_q , \slAcky/mxl/muxout , \slAckx/l1_q , 
        \slAckx/mxl/muxout ;
    nor2_2 U12 ( .x(nack_x), .a(ackx_l), .b(rst) );
    nand2_1 U4 ( .x(ack_ix), .a(n1x), .b(n2x) );
    nor3_1 U17 ( .x(n1x), .a(d2_ox), .b(d3_ox), .c(d1_ox) );
    nor2_1 U18 ( .x(n2x), .a(eop_ox), .b(d0_ox) );
    nor2_2 U11 ( .x(nack_y), .a(acky_l), .b(rst) );
    nand2_1 U3 ( .x(ack_iy), .a(n1y), .b(n2y) );
    nor3_1 U16 ( .x(n1y), .a(d2_oy), .b(d3_oy), .c(d1_oy) );
    nor2_1 U19 ( .x(n2y), .a(eop_oy), .b(d0_oy) );
    nand2_1 U15 ( .x(req_x), .a(n5x), .b(n6x) );
    nor3_1 U10 ( .x(n5x), .a(d2_ix), .b(d3_ix), .c(d1_ix) );
    nor2_1 U13 ( .x(n6x), .a(eop_ix), .b(d0_ix) );
    nand2_1 U14 ( .x(req_y), .a(n5y), .b(n6y) );
    nor3_1 U9 ( .x(n5y), .a(d2_iy), .b(d3_iy), .c(d1_iy) );
    nor2_1 U20 ( .x(n6y), .a(eop_iy), .b(d0_iy) );
    nor2i_1 U6 ( .x(sx_pl), .a(gx), .b(eop_oy) );
    nor2i_1 U5 ( .x(sy_pl), .a(gy), .b(eop_ox) );
    nor3_1 \cye/Unr  ( .x(\cye/nr ), .a(eop_iy), .b(nack_y), .c(sy) );
    nand3_1 \cye/Und  ( .x(\cye/nd ), .a(eop_iy), .b(nack_y), .c(sy) );
    oa21_1 \cye/U1  ( .x(\cye/n2 ), .a(\cye/n2 ), .b(\cye/nr ), .c(\cye/nd )
         );
    inv_1 \cye/U3  ( .x(eop_oy), .a(\cye/n2 ) );
    ao31_1 \cy3/__tmp99/aoi  ( .x(\cy3/__tmp99/loop ), .a(d3_iy), .b(nack_y), 
        .c(sy), .d(d3_oy) );
    oa21_1 \cy3/__tmp99/outGate  ( .x(d3_oy), .a(d3_iy), .b(nack_y), .c(
        \cy3/__tmp99/loop ) );
    ao31_1 \cy2/__tmp99/aoi  ( .x(\cy2/__tmp99/loop ), .a(d2_iy), .b(nack_y), 
        .c(sy), .d(d2_oy) );
    oa21_1 \cy2/__tmp99/outGate  ( .x(d2_oy), .a(d2_iy), .b(nack_y), .c(
        \cy2/__tmp99/loop ) );
    ao31_1 \cy1/__tmp99/aoi  ( .x(\cy1/__tmp99/loop ), .a(d1_iy), .b(nack_y), 
        .c(sy), .d(d1_oy) );
    oa21_1 \cy1/__tmp99/outGate  ( .x(d1_oy), .a(d1_iy), .b(nack_y), .c(
        \cy1/__tmp99/loop ) );
    ao31_1 \cy0/__tmp99/aoi  ( .x(\cy0/__tmp99/loop ), .a(d0_iy), .b(nack_y), 
        .c(sy), .d(d0_oy) );
    oa21_1 \cy0/__tmp99/outGate  ( .x(d0_oy), .a(d0_iy), .b(nack_y), .c(
        \cy0/__tmp99/loop ) );
    nor3_1 \cxe/Unr  ( .x(\cxe/nr ), .a(eop_ix), .b(nack_x), .c(sx) );
    nand3_1 \cxe/Und  ( .x(\cxe/nd ), .a(eop_ix), .b(nack_x), .c(sx) );
    oa21_1 \cxe/U1  ( .x(\cxe/n2 ), .a(\cxe/n2 ), .b(\cxe/nr ), .c(\cxe/nd )
         );
    inv_1 \cxe/U3  ( .x(eop_ox), .a(\cxe/n2 ) );
    ao31_1 \cx3/__tmp99/aoi  ( .x(\cx3/__tmp99/loop ), .a(d3_ix), .b(nack_x), 
        .c(sx), .d(d3_ox) );
    oa21_1 \cx3/__tmp99/outGate  ( .x(d3_ox), .a(d3_ix), .b(nack_x), .c(
        \cx3/__tmp99/loop ) );
    ao31_1 \cx2/__tmp99/aoi  ( .x(\cx2/__tmp99/loop ), .a(d2_ix), .b(nack_x), 
        .c(sx), .d(d2_ox) );
    oa21_1 \cx2/__tmp99/outGate  ( .x(d2_ox), .a(d2_ix), .b(nack_x), .c(
        \cx2/__tmp99/loop ) );
    ao31_1 \cx1/__tmp99/aoi  ( .x(\cx1/__tmp99/loop ), .a(d1_ix), .b(nack_x), 
        .c(sx), .d(d1_ox) );
    oa21_1 \cx1/__tmp99/outGate  ( .x(d1_ox), .a(d1_ix), .b(nack_x), .c(
        \cx1/__tmp99/loop ) );
    ao31_1 \cx0/__tmp99/aoi  ( .x(\cx0/__tmp99/loop ), .a(d0_ix), .b(nack_x), 
        .c(sx), .d(d0_ox) );
    oa21_1 \cx0/__tmp99/outGate  ( .x(d0_ox), .a(d0_ix), .b(nack_x), .c(
        \cx0/__tmp99/loop ) );
    nand2_1 \mtx/mg2  ( .x(\mtx/gr2 ), .a(mry), .b(\mtx/gr1 ) );
    nand2_1 \mtx/U1  ( .x(\mtx/gr1 ), .a(mrx), .b(\mtx/gr2 ) );
    nor3_1 \mtx/U2  ( .x(gy), .a(\mtx/gr2 ), .b(\mtx/gr2 ), .c(\mtx/gr2 ) );
    nor3_1 \mtx/U3  ( .x(gx), .a(\mtx/gr1 ), .b(\mtx/gr1 ), .c(\mtx/gr1 ) );
    nor2_1 \sry/i1  ( .x(\sry/qz ), .a(req_y), .b(mry) );
    nor2_1 \srx/i1  ( .x(\srx/qz ), .a(req_x), .b(mrx) );
    latn_1 \sl_sy/lph3  ( .q(sy), .d(\sl_sy/l1_q ), .g(phi3) );
    latn_1 \sl_sy/lph2  ( .q(\scan[1] ), .d(\sl_sy/l1_q ), .g(phi2) );
    mux2_1 \sl_sy/mxl/mux  ( .x(\sl_sy/mxl/muxout ), .d0(sy_pl), .sl(test_se), 
        .d1(\scan[0] ) );
    latn_1 \sl_sy/mxl/lph1  ( .q(\sl_sy/l1_q ), .d(\sl_sy/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_sx/lph3  ( .q(sx), .d(\sl_sx/l1_q ), .g(phi3) );
    latn_1 \sl_sx/lph2  ( .q(\scan[0] ), .d(\sl_sx/l1_q ), .g(phi2) );
    mux2_1 \sl_sx/mxl/mux  ( .x(\sl_sx/mxl/muxout ), .d0(sx_pl), .sl(test_se), 
        .d1(test_si) );
    latn_1 \sl_sx/mxl/lph1  ( .q(\sl_sx/l1_q ), .d(\sl_sx/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAcky/lph3  ( .q(acky_l), .d(\slAcky/l1_q ), .g(phi3) );
    latn_1 \slAcky/lph2  ( .q(test_so), .d(\slAcky/l1_q ), .g(phi2) );
    mux2_1 \slAcky/mxl/mux  ( .x(\slAcky/mxl/muxout ), .d0(ack_oxy), .sl(
        test_se), .d1(\scan[2] ) );
    latn_1 \slAcky/mxl/lph1  ( .q(\slAcky/l1_q ), .d(\slAcky/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAckx/lph3  ( .q(ackx_l), .d(\slAckx/l1_q ), .g(phi3) );
    latn_1 \slAckx/lph2  ( .q(\scan[2] ), .d(\slAckx/l1_q ), .g(phi2) );
    mux2_1 \slAckx/mxl/mux  ( .x(\slAckx/mxl/muxout ), .d0(ack_oxy), .sl(
        test_se), .d1(\scan[1] ) );
    latn_1 \slAckx/mxl/lph1  ( .q(\slAckx/l1_q ), .d(\slAckx/mxl/muxout ), .g(
        phi1) );
    nor3_0 U1 ( .x(mrx), .a(eop_ox), .b(rst), .c(\srx/qz ) );
    nor3_1 U2 ( .x(mry), .a(eop_oy), .b(rst), .c(\sry/qz ) );
endmodule


module chain_arbiter1 ( eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, ack_ix, eop_iy, 
    d0_iy, d1_iy, d2_iy, d3_iy, ack_iy, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, 
    eop_oy, d0_oy, d1_oy, d2_oy, d3_oy, ack_oxy, rst, test_si, test_se, 
    test_so, phi1, phi2, phi3 );
input  eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, eop_iy, d0_iy, d1_iy, d2_iy, d3_iy, 
    ack_oxy, rst, test_si, test_se, phi1, phi2, phi3;
output ack_ix, ack_iy, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, eop_oy, d0_oy, 
    d1_oy, d2_oy, d3_oy, test_so;
    wire \scan[1] , \scan[2] , ackx_l, nack_x, sx, acky_l, nack_y, sy, mrx, 
        req_x, mry, req_y, gx, gy, \scan[0] , sx_pl, sy_pl, n1x, n2x, n1y, n2y, 
        n5x, n6x, n5y, n6y, \cye/nr , \cye/nd , \cye/n2 , \cy3/__tmp99/loop , 
        \cy2/__tmp99/loop , \cy1/__tmp99/loop , \cy0/__tmp99/loop , \cxe/nr , 
        \cxe/nd , \cxe/n2 , \cx3/__tmp99/loop , \cx2/__tmp99/loop , 
        \cx1/__tmp99/loop , \cx0/__tmp99/loop , \mtx/gr2 , \mtx/gr1 , \sry/qz , 
        \srx/qz , \sl_sy/l1_q , \sl_sy/mxl/muxout , \sl_sx/l1_q , 
        \sl_sx/mxl/muxout , \slAcky/l1_q , \slAcky/mxl/muxout , \slAckx/l1_q , 
        \slAckx/mxl/muxout ;
    nor2_2 U12 ( .x(nack_x), .a(ackx_l), .b(rst) );
    nand2_1 U4 ( .x(ack_ix), .a(n1x), .b(n2x) );
    nor3_1 U17 ( .x(n1x), .a(d2_ox), .b(d3_ox), .c(d1_ox) );
    nor2_1 U18 ( .x(n2x), .a(eop_ox), .b(d0_ox) );
    nor2_2 U11 ( .x(nack_y), .a(acky_l), .b(rst) );
    nand2_1 U3 ( .x(ack_iy), .a(n1y), .b(n2y) );
    nor3_1 U16 ( .x(n1y), .a(d2_oy), .b(d3_oy), .c(d1_oy) );
    nor2_1 U19 ( .x(n2y), .a(eop_oy), .b(d0_oy) );
    nand2_1 U15 ( .x(req_x), .a(n5x), .b(n6x) );
    nor3_1 U10 ( .x(n5x), .a(d2_ix), .b(d3_ix), .c(d1_ix) );
    nor2_1 U13 ( .x(n6x), .a(eop_ix), .b(d0_ix) );
    nand2_1 U14 ( .x(req_y), .a(n5y), .b(n6y) );
    nor3_1 U9 ( .x(n5y), .a(d2_iy), .b(d3_iy), .c(d1_iy) );
    nor2_1 U20 ( .x(n6y), .a(eop_iy), .b(d0_iy) );
    nor2i_1 U6 ( .x(sx_pl), .a(gx), .b(eop_oy) );
    nor2i_1 U5 ( .x(sy_pl), .a(gy), .b(eop_ox) );
    nor3_1 \cye/Unr  ( .x(\cye/nr ), .a(eop_iy), .b(nack_y), .c(sy) );
    nand3_1 \cye/Und  ( .x(\cye/nd ), .a(eop_iy), .b(nack_y), .c(sy) );
    oa21_1 \cye/U1  ( .x(\cye/n2 ), .a(\cye/n2 ), .b(\cye/nr ), .c(\cye/nd )
         );
    inv_1 \cye/U3  ( .x(eop_oy), .a(\cye/n2 ) );
    ao31_1 \cy3/__tmp99/aoi  ( .x(\cy3/__tmp99/loop ), .a(d3_iy), .b(nack_y), 
        .c(sy), .d(d3_oy) );
    oa21_1 \cy3/__tmp99/outGate  ( .x(d3_oy), .a(d3_iy), .b(nack_y), .c(
        \cy3/__tmp99/loop ) );
    ao31_1 \cy2/__tmp99/aoi  ( .x(\cy2/__tmp99/loop ), .a(d2_iy), .b(nack_y), 
        .c(sy), .d(d2_oy) );
    oa21_1 \cy2/__tmp99/outGate  ( .x(d2_oy), .a(d2_iy), .b(nack_y), .c(
        \cy2/__tmp99/loop ) );
    ao31_1 \cy1/__tmp99/aoi  ( .x(\cy1/__tmp99/loop ), .a(d1_iy), .b(nack_y), 
        .c(sy), .d(d1_oy) );
    oa21_1 \cy1/__tmp99/outGate  ( .x(d1_oy), .a(d1_iy), .b(nack_y), .c(
        \cy1/__tmp99/loop ) );
    ao31_1 \cy0/__tmp99/aoi  ( .x(\cy0/__tmp99/loop ), .a(d0_iy), .b(nack_y), 
        .c(sy), .d(d0_oy) );
    oa21_1 \cy0/__tmp99/outGate  ( .x(d0_oy), .a(d0_iy), .b(nack_y), .c(
        \cy0/__tmp99/loop ) );
    nor3_1 \cxe/Unr  ( .x(\cxe/nr ), .a(eop_ix), .b(nack_x), .c(sx) );
    nand3_1 \cxe/Und  ( .x(\cxe/nd ), .a(eop_ix), .b(nack_x), .c(sx) );
    oa21_1 \cxe/U1  ( .x(\cxe/n2 ), .a(\cxe/n2 ), .b(\cxe/nr ), .c(\cxe/nd )
         );
    inv_1 \cxe/U3  ( .x(eop_ox), .a(\cxe/n2 ) );
    ao31_1 \cx3/__tmp99/aoi  ( .x(\cx3/__tmp99/loop ), .a(d3_ix), .b(nack_x), 
        .c(sx), .d(d3_ox) );
    oa21_1 \cx3/__tmp99/outGate  ( .x(d3_ox), .a(d3_ix), .b(nack_x), .c(
        \cx3/__tmp99/loop ) );
    ao31_1 \cx2/__tmp99/aoi  ( .x(\cx2/__tmp99/loop ), .a(d2_ix), .b(nack_x), 
        .c(sx), .d(d2_ox) );
    oa21_1 \cx2/__tmp99/outGate  ( .x(d2_ox), .a(d2_ix), .b(nack_x), .c(
        \cx2/__tmp99/loop ) );
    ao31_1 \cx1/__tmp99/aoi  ( .x(\cx1/__tmp99/loop ), .a(d1_ix), .b(nack_x), 
        .c(sx), .d(d1_ox) );
    oa21_1 \cx1/__tmp99/outGate  ( .x(d1_ox), .a(d1_ix), .b(nack_x), .c(
        \cx1/__tmp99/loop ) );
    ao31_1 \cx0/__tmp99/aoi  ( .x(\cx0/__tmp99/loop ), .a(d0_ix), .b(nack_x), 
        .c(sx), .d(d0_ox) );
    oa21_1 \cx0/__tmp99/outGate  ( .x(d0_ox), .a(d0_ix), .b(nack_x), .c(
        \cx0/__tmp99/loop ) );
    nand2_1 \mtx/mg2  ( .x(\mtx/gr2 ), .a(mry), .b(\mtx/gr1 ) );
    nand2_1 \mtx/U1  ( .x(\mtx/gr1 ), .a(mrx), .b(\mtx/gr2 ) );
    nor3_1 \mtx/U2  ( .x(gy), .a(\mtx/gr2 ), .b(\mtx/gr2 ), .c(\mtx/gr2 ) );
    nor3_1 \mtx/U3  ( .x(gx), .a(\mtx/gr1 ), .b(\mtx/gr1 ), .c(\mtx/gr1 ) );
    nor2_1 \sry/i1  ( .x(\sry/qz ), .a(req_y), .b(mry) );
    nor2_1 \srx/i1  ( .x(\srx/qz ), .a(req_x), .b(mrx) );
    latn_1 \sl_sy/lph3  ( .q(sy), .d(\sl_sy/l1_q ), .g(phi3) );
    latn_1 \sl_sy/lph2  ( .q(\scan[1] ), .d(\sl_sy/l1_q ), .g(phi2) );
    mux2_1 \sl_sy/mxl/mux  ( .x(\sl_sy/mxl/muxout ), .d0(sy_pl), .sl(test_se), 
        .d1(\scan[0] ) );
    latn_1 \sl_sy/mxl/lph1  ( .q(\sl_sy/l1_q ), .d(\sl_sy/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_sx/lph3  ( .q(sx), .d(\sl_sx/l1_q ), .g(phi3) );
    latn_1 \sl_sx/lph2  ( .q(\scan[0] ), .d(\sl_sx/l1_q ), .g(phi2) );
    mux2_1 \sl_sx/mxl/mux  ( .x(\sl_sx/mxl/muxout ), .d0(sx_pl), .sl(test_se), 
        .d1(test_si) );
    latn_1 \sl_sx/mxl/lph1  ( .q(\sl_sx/l1_q ), .d(\sl_sx/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAcky/lph3  ( .q(acky_l), .d(\slAcky/l1_q ), .g(phi3) );
    latn_1 \slAcky/lph2  ( .q(test_so), .d(\slAcky/l1_q ), .g(phi2) );
    mux2_1 \slAcky/mxl/mux  ( .x(\slAcky/mxl/muxout ), .d0(ack_oxy), .sl(
        test_se), .d1(\scan[2] ) );
    latn_1 \slAcky/mxl/lph1  ( .q(\slAcky/l1_q ), .d(\slAcky/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAckx/lph3  ( .q(ackx_l), .d(\slAckx/l1_q ), .g(phi3) );
    latn_1 \slAckx/lph2  ( .q(\scan[2] ), .d(\slAckx/l1_q ), .g(phi2) );
    mux2_1 \slAckx/mxl/mux  ( .x(\slAckx/mxl/muxout ), .d0(ack_oxy), .sl(
        test_se), .d1(\scan[1] ) );
    latn_1 \slAckx/mxl/lph1  ( .q(\slAckx/l1_q ), .d(\slAckx/mxl/muxout ), .g(
        phi1) );
    nor3_1 U1 ( .x(mrx), .a(eop_ox), .b(rst), .c(\srx/qz ) );
    nor3_1 U2 ( .x(mry), .a(eop_oy), .b(rst), .c(\sry/qz ) );
endmodule


module chain_mux0 ( eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, ack_ixy, eop_iy, d0_iy, 
    d1_iy, d2_iy, d3_iy, eop_o, d0_o, d1_o, d2_o, d3_o, ack_o, rst, test_si, 
    test_se, test_so, phi1, phi2, phi3 );
input  eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, eop_iy, d0_iy, d1_iy, d2_iy, d3_iy, 
    ack_o, rst, test_si, test_se, phi1, phi2, phi3;
output ack_ixy, eop_o, d0_o, d1_o, d2_o, d3_o, test_so;
    wire ack_l, d0_i, ack, d1_i, d2_i, d3_i, eop_i, n1, n2, \ce/ob , \c3/ob , 
        \c2/ob , \c1/ob , \c0/ob , \slAck/l1_q , \slAck/mxl/muxout ;
    nor2_1 U2 ( .x(d3_i), .a(d3_iy), .b(d3_ix) );
    nor2_1 U3 ( .x(d2_i), .a(d2_iy), .b(d2_ix) );
    nor2_1 U4 ( .x(d1_i), .a(d1_iy), .b(d1_ix) );
    nor2_1 U5 ( .x(d0_i), .a(d0_iy), .b(d0_ix) );
    nor2_1 U6 ( .x(eop_i), .a(eop_iy), .b(eop_ix) );
    nand2_1 U1 ( .x(ack_ixy), .a(n1), .b(n2) );
    nor3_1 U9 ( .x(n1), .a(d2_o), .b(d3_o), .c(d1_o) );
    nor2_1 U8 ( .x(n2), .a(eop_o), .b(d0_o) );
    inv_1 \ce/Ui  ( .x(\ce/ob ), .a(eop_o) );
    aoi222_1 \ce/__tmp99/U1  ( .x(eop_o), .a(eop_i), .b(ack), .c(eop_i), .d(
        \ce/ob ), .e(ack), .f(\ce/ob ) );
    inv_1 \c3/Ui  ( .x(\c3/ob ), .a(d3_o) );
    aoi222_1 \c3/__tmp99/U1  ( .x(d3_o), .a(d3_i), .b(ack), .c(d3_i), .d(
        \c3/ob ), .e(ack), .f(\c3/ob ) );
    inv_1 \c2/Ui  ( .x(\c2/ob ), .a(d2_o) );
    aoi222_1 \c2/__tmp99/U1  ( .x(d2_o), .a(d2_i), .b(ack), .c(d2_i), .d(
        \c2/ob ), .e(ack), .f(\c2/ob ) );
    inv_1 \c1/Ui  ( .x(\c1/ob ), .a(d1_o) );
    aoi222_1 \c1/__tmp99/U1  ( .x(d1_o), .a(d1_i), .b(ack), .c(d1_i), .d(
        \c1/ob ), .e(ack), .f(\c1/ob ) );
    inv_1 \c0/Ui  ( .x(\c0/ob ), .a(d0_o) );
    aoi222_1 \c0/__tmp99/U1  ( .x(d0_o), .a(d0_i), .b(ack), .c(d0_i), .d(
        \c0/ob ), .e(ack), .f(\c0/ob ) );
    latn_1 \slAck/lph3  ( .q(ack_l), .d(\slAck/l1_q ), .g(phi3) );
    latn_1 \slAck/lph2  ( .q(test_so), .d(\slAck/l1_q ), .g(phi2) );
    mux2_1 \slAck/mxl/mux  ( .x(\slAck/mxl/muxout ), .d0(ack_o), .sl(test_se), 
        .d1(test_si) );
    latn_1 \slAck/mxl/lph1  ( .q(\slAck/l1_q ), .d(\slAck/mxl/muxout ), .g(
        phi1) );
    or2_3 U7 ( .x(ack), .a(ack_l), .b(rst) );
endmodule


module chain_mux1 ( eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, ack_ixy, eop_iy, d0_iy, 
    d1_iy, d2_iy, d3_iy, eop_o, d0_o, d1_o, d2_o, d3_o, ack_o, rst, test_si, 
    test_se, test_so, phi1, phi2, phi3 );
input  eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, eop_iy, d0_iy, d1_iy, d2_iy, d3_iy, 
    ack_o, rst, test_si, test_se, phi1, phi2, phi3;
output ack_ixy, eop_o, d0_o, d1_o, d2_o, d3_o, test_so;
    wire ack_l, d0_i, ack, d1_i, d2_i, d3_i, eop_i, n1, n2, \ce/ob , \c3/ob , 
        \c2/ob , \c1/ob , \c0/ob , \slAck/l1_q , \slAck/mxl/muxout ;
    nor2_1 U2 ( .x(d3_i), .a(d3_iy), .b(d3_ix) );
    nor2_1 U3 ( .x(d2_i), .a(d2_iy), .b(d2_ix) );
    nor2_1 U4 ( .x(d1_i), .a(d1_iy), .b(d1_ix) );
    nor2_1 U5 ( .x(d0_i), .a(d0_iy), .b(d0_ix) );
    nor2_1 U6 ( .x(eop_i), .a(eop_iy), .b(eop_ix) );
    nand2_1 U1 ( .x(ack_ixy), .a(n1), .b(n2) );
    nor3_1 U9 ( .x(n1), .a(d2_o), .b(d3_o), .c(d1_o) );
    nor2_1 U8 ( .x(n2), .a(eop_o), .b(d0_o) );
    inv_1 \ce/Ui  ( .x(\ce/ob ), .a(eop_o) );
    aoi222_1 \ce/__tmp99/U1  ( .x(eop_o), .a(eop_i), .b(ack), .c(eop_i), .d(
        \ce/ob ), .e(ack), .f(\ce/ob ) );
    inv_1 \c3/Ui  ( .x(\c3/ob ), .a(d3_o) );
    aoi222_1 \c3/__tmp99/U1  ( .x(d3_o), .a(d3_i), .b(ack), .c(d3_i), .d(
        \c3/ob ), .e(ack), .f(\c3/ob ) );
    inv_1 \c2/Ui  ( .x(\c2/ob ), .a(d2_o) );
    aoi222_1 \c2/__tmp99/U1  ( .x(d2_o), .a(d2_i), .b(ack), .c(d2_i), .d(
        \c2/ob ), .e(ack), .f(\c2/ob ) );
    inv_1 \c1/Ui  ( .x(\c1/ob ), .a(d1_o) );
    aoi222_1 \c1/__tmp99/U1  ( .x(d1_o), .a(d1_i), .b(ack), .c(d1_i), .d(
        \c1/ob ), .e(ack), .f(\c1/ob ) );
    inv_1 \c0/Ui  ( .x(\c0/ob ), .a(d0_o) );
    aoi222_1 \c0/__tmp99/U1  ( .x(d0_o), .a(d0_i), .b(ack), .c(d0_i), .d(
        \c0/ob ), .e(ack), .f(\c0/ob ) );
    latn_1 \slAck/lph3  ( .q(ack_l), .d(\slAck/l1_q ), .g(phi3) );
    latn_1 \slAck/lph2  ( .q(test_so), .d(\slAck/l1_q ), .g(phi2) );
    mux2_1 \slAck/mxl/mux  ( .x(\slAck/mxl/muxout ), .d0(ack_o), .sl(test_se), 
        .d1(test_si) );
    latn_1 \slAck/mxl/lph1  ( .q(\slAck/l1_q ), .d(\slAck/mxl/muxout ), .g(
        phi1) );
    or2_3 U7 ( .x(ack), .a(ack_l), .b(rst) );
endmodule


module comm_fab ( nrst, I_port_eop_i, I_port_d0_i, I_port_d1_i, I_port_d2_i, 
    I_port_d3_i, I_port_ack, TIC_eop_i, TIC_d0_i, TIC_d1_i, TIC_d2_i, TIC_d3_i, 
    TIC_ack, D_port_eop_i, D_port_d0_i, D_port_d1_i, D_port_d2_i, D_port_d3_i, 
    D_port_ack, BC_eop_i, BC_d0_i, BC_d1_i, BC_d2_i, BC_d3_i, BC_ack, WB_eop_i, 
    WB_d0_i, WB_d1_i, WB_d2_i, WB_d3_i, WB_ack, IMEM_eop_i, IMEM_d0_i, 
    IMEM_d1_i, IMEM_d2_i, IMEM_d3_i, IMEM_ack, DMEM_eop_i, DMEM_d0_i, 
    DMEM_d1_i, DMEM_d2_i, DMEM_d3_i, DMEM_ack, test_si, test_so, test_se, phi1, 
    phi2, phi3 );
input  nrst, I_port_eop_i, I_port_d0_i, I_port_d1_i, I_port_d2_i, I_port_d3_i, 
    TIC_eop_i, TIC_d0_i, TIC_d1_i, TIC_d2_i, TIC_d3_i, D_port_eop_i, 
    D_port_d0_i, D_port_d1_i, D_port_d2_i, D_port_d3_i, BC_ack, WB_ack, 
    IMEM_ack, DMEM_ack, test_si, test_se, phi1, phi2, phi3;
output I_port_ack, TIC_ack, D_port_ack, BC_eop_i, BC_d0_i, BC_d1_i, BC_d2_i, 
    BC_d3_i, WB_eop_i, WB_d0_i, WB_d1_i, WB_d2_i, WB_d3_i, IMEM_eop_i, 
    IMEM_d0_i, IMEM_d1_i, IMEM_d2_i, IMEM_d3_i, DMEM_eop_i, DMEM_d0_i, 
    DMEM_d1_i, DMEM_d2_i, DMEM_d3_i, test_so;
    wire rst, A0_eop_o0, A0_d0_o0, A0_d1_o0, A0_d2_o0, A0_d3_o0, A0_eop_o1, 
        A0_d0_o1, A0_d1_o1, A0_d2_o1, A0_d3_o1, A0_ack, \scan[6] , \scan[5] , 
        \scan[4] , \scan[3] , \scan[2] , \scan[1] , M0_eop, M0_d0, M0_d1, 
        M0_d2, M0_d3, M0_ack, A1_eop_o0, A1_d0_o0, A1_d1_o0, A1_d2_o0, 
        A1_d3_o0, A1_eop_o1, A1_d0_o1, A1_d1_o1, A1_d2_o1, A1_d3_o1, A1_ack, 
        M1_eop, M1_d0, M1_d1, M1_d2, M1_d3, M1_ack, R0_odd_eop, R0_odd_d0, 
        R0_odd_d1, R0_odd_d2, R0_odd_d3, R0_odd_ack, R1_odd_eop, R1_odd_d0, 
        R1_odd_d1, R1_odd_d2, R1_odd_d3, R1_odd_ack, n1, n2, n3, n4;
    inv_2 U1 ( .x(rst), .a(nrst) );
    chain_arbiter0 arb0 ( .eop_ix(I_port_eop_i), .d0_ix(I_port_d0_i), .d1_ix(
        I_port_d1_i), .d2_ix(I_port_d2_i), .d3_ix(I_port_d3_i), .ack_ix(
        I_port_ack), .eop_iy(D_port_eop_i), .d0_iy(D_port_d0_i), .d1_iy(
        D_port_d1_i), .d2_iy(D_port_d2_i), .d3_iy(D_port_d3_i), .ack_iy(
        D_port_ack), .eop_ox(A0_eop_o0), .d0_ox(A0_d0_o0), .d1_ox(A0_d1_o0), 
        .d2_ox(A0_d2_o0), .d3_ox(A0_d3_o0), .eop_oy(A0_eop_o1), .d0_oy(
        A0_d0_o1), .d1_oy(A0_d1_o1), .d2_oy(A0_d2_o1), .d3_oy(A0_d3_o1), 
        .ack_oxy(A0_ack), .rst(rst), .test_si(test_si), .test_se(n4), 
        .test_so(\scan[1] ), .phi1(phi1), .phi2(phi2), .phi3(phi3) );
    chain_mux0 mux0 ( .eop_ix(A0_eop_o0), .d0_ix(A0_d0_o0), .d1_ix(A0_d1_o0), 
        .d2_ix(A0_d2_o0), .d3_ix(A0_d3_o0), .ack_ixy(A0_ack), .eop_iy(
        A0_eop_o1), .d0_iy(A0_d0_o1), .d1_iy(A0_d1_o1), .d2_iy(A0_d2_o1), 
        .d3_iy(A0_d3_o1), .eop_o(M0_eop), .d0_o(M0_d0), .d1_o(M0_d1), .d2_o(
        M0_d2), .d3_o(M0_d3), .ack_o(M0_ack), .rst(rst), .test_si(\scan[1] ), 
        .test_se(n4), .test_so(\scan[2] ), .phi1(n2), .phi2(n1), .phi3(n3) );
    chain_arbiter1 arb1 ( .eop_ix(M0_eop), .d0_ix(M0_d0), .d1_ix(M0_d1), 
        .d2_ix(M0_d2), .d3_ix(M0_d3), .ack_ix(M0_ack), .eop_iy(TIC_eop_i), 
        .d0_iy(TIC_d0_i), .d1_iy(TIC_d1_i), .d2_iy(TIC_d2_i), .d3_iy(TIC_d3_i), 
        .ack_iy(TIC_ack), .eop_ox(A1_eop_o0), .d0_ox(A1_d0_o0), .d1_ox(
        A1_d1_o0), .d2_ox(A1_d2_o0), .d3_ox(A1_d3_o0), .eop_oy(A1_eop_o1), 
        .d0_oy(A1_d0_o1), .d1_oy(A1_d1_o1), .d2_oy(A1_d2_o1), .d3_oy(A1_d3_o1), 
        .ack_oxy(A1_ack), .rst(rst), .test_si(\scan[2] ), .test_se(n4), 
        .test_so(\scan[3] ), .phi1(n2), .phi2(n1), .phi3(n3) );
    chain_mux1 mux1 ( .eop_ix(A1_eop_o0), .d0_ix(A1_d0_o0), .d1_ix(A1_d1_o0), 
        .d2_ix(A1_d2_o0), .d3_ix(A1_d3_o0), .ack_ixy(A1_ack), .eop_iy(
        A1_eop_o1), .d0_iy(A1_d0_o1), .d1_iy(A1_d1_o1), .d2_iy(A1_d2_o1), 
        .d3_iy(A1_d3_o1), .eop_o(M1_eop), .d0_o(M1_d0), .d1_o(M1_d1), .d2_o(
        M1_d2), .d3_o(M1_d3), .ack_o(M1_ack), .rst(rst), .test_si(\scan[3] ), 
        .test_se(test_se), .test_so(\scan[4] ), .phi1(phi1), .phi2(phi2), 
        .phi3(phi3) );
    chain_router0 router0 ( .eop_i(M1_eop), .d0_i(M1_d0), .d1_i(M1_d1), .d2_i(
        M1_d2), .d3_i(M1_d3), .ack_i(M1_ack), .eop_ox(R0_odd_eop), .d0_ox(
        R0_odd_d0), .d1_ox(R0_odd_d1), .d2_ox(R0_odd_d2), .d3_ox(R0_odd_d3), 
        .ack_ox(R0_odd_ack), .eop_oy(WB_eop_i), .d0_oy(WB_d0_i), .d1_oy(
        WB_d1_i), .d2_oy(WB_d2_i), .d3_oy(WB_d3_i), .ack_oy(WB_ack), .nrst(
        nrst), .test_si(\scan[4] ), .test_se(test_se), .test_so(\scan[5] ), 
        .phi1(phi1), .phi2(phi2), .phi3(phi3) );
    chain_router1 router1 ( .eop_i(R0_odd_eop), .d0_i(R0_odd_d0), .d1_i(
        R0_odd_d1), .d2_i(R0_odd_d2), .d3_i(R0_odd_d3), .ack_i(R0_odd_ack), 
        .eop_ox(R1_odd_eop), .d0_ox(R1_odd_d0), .d1_ox(R1_odd_d1), .d2_ox(
        R1_odd_d2), .d3_ox(R1_odd_d3), .ack_ox(R1_odd_ack), .eop_oy(BC_eop_i), 
        .d0_oy(BC_d0_i), .d1_oy(BC_d1_i), .d2_oy(BC_d2_i), .d3_oy(BC_d3_i), 
        .ack_oy(BC_ack), .nrst(nrst), .test_si(\scan[5] ), .test_se(n4), 
        .test_so(\scan[6] ), .phi1(n2), .phi2(n1), .phi3(n3) );
    chain_router2 router2 ( .eop_i(R1_odd_eop), .d0_i(R1_odd_d0), .d1_i(
        R1_odd_d1), .d2_i(R1_odd_d2), .d3_i(R1_odd_d3), .ack_i(R1_odd_ack), 
        .eop_ox(DMEM_eop_i), .d0_ox(DMEM_d0_i), .d1_ox(DMEM_d1_i), .d2_ox(
        DMEM_d2_i), .d3_ox(DMEM_d3_i), .ack_ox(DMEM_ack), .eop_oy(IMEM_eop_i), 
        .d0_oy(IMEM_d0_i), .d1_oy(IMEM_d1_i), .d2_oy(IMEM_d2_i), .d3_oy(
        IMEM_d3_i), .ack_oy(IMEM_ack), .nrst(nrst), .test_si(\scan[6] ), 
        .test_se(test_se), .test_so(test_so), .phi1(phi1), .phi2(phi2), .phi3(
        phi3) );
    buf_1 U2 ( .x(n1), .a(phi2) );
    buf_1 U3 ( .x(n2), .a(phi1) );
    buf_1 U4 ( .x(n3), .a(phi3) );
    buf_3 U5 ( .x(n4), .a(test_se) );
endmodule


module comm_fab_scan ( nrst, I_port_eop_i, I_port_d0_i, I_port_d1_i, 
    I_port_d2_i, I_port_d3_i, I_port_ack, TIC_eop_i, TIC_d0_i, TIC_d1_i, 
    TIC_d2_i, TIC_d3_i, TIC_ack, D_port_eop_i, D_port_d0_i, D_port_d1_i, 
    D_port_d2_i, D_port_d3_i, D_port_ack, BC_eop_i, BC_d0_i, BC_d1_i, BC_d2_i, 
    BC_d3_i, BC_ack, WB_eop_i, WB_d0_i, WB_d1_i, WB_d2_i, WB_d3_i, WB_ack, 
    IMEM_eop_i, IMEM_d0_i, IMEM_d1_i, IMEM_d2_i, IMEM_d3_i, IMEM_ack, 
    DMEM_eop_i, DMEM_d0_i, DMEM_d1_i, DMEM_d2_i, DMEM_d3_i, DMEM_ack, test_si, 
    test_so, test_se, phi1, phi2, phi3 );
input  nrst, I_port_eop_i, I_port_d0_i, I_port_d1_i, I_port_d2_i, I_port_d3_i, 
    TIC_eop_i, TIC_d0_i, TIC_d1_i, TIC_d2_i, TIC_d3_i, D_port_eop_i, 
    D_port_d0_i, D_port_d1_i, D_port_d2_i, D_port_d3_i, BC_ack, WB_ack, 
    IMEM_ack, DMEM_ack, test_si, test_se, phi1, phi2, phi3;
output I_port_ack, TIC_ack, D_port_ack, BC_eop_i, BC_d0_i, BC_d1_i, BC_d2_i, 
    BC_d3_i, WB_eop_i, WB_d0_i, WB_d1_i, WB_d2_i, WB_d3_i, IMEM_eop_i, 
    IMEM_d0_i, IMEM_d1_i, IMEM_d2_i, IMEM_d3_i, DMEM_eop_i, DMEM_d0_i, 
    DMEM_d1_i, DMEM_d2_i, DMEM_d3_i, test_so;
    wire \scan[12] , \scan[11] , \scan[10] , \scan[9] , \scan[8] , \scan[7] , 
        \scan[6] , \scan[5] , \scan[4] , \scan[3] , \scan[2] , \scan[1] , 
        I_port_eop_i_sc, I_port_d0_i_sc, I_port_d1_i_sc, I_port_d2_i_sc, 
        I_port_d3_i_sc, TIC_eop_i_sc, TIC_d0_i_sc, TIC_d1_i_sc, TIC_d2_i_sc, 
        TIC_d3_i_sc, D_port_eop_i_sc, D_port_d0_i_sc, D_port_d1_i_sc, 
        D_port_d2_i_sc, D_port_d3_i_sc, WB_ack_sc, IMEM_ack_sc, DMEM_ack_sc, 
        scan_m10, scan_m11, scan_m12, \sc12_m_dpAck/muxout , 
        \sc11_m_ticAck/muxout , \sc10_m_ipAck/muxout , \sc5_dmAck/l1_q , 
        \sc5_dmAck/mxl/muxout , \sc4_imAck/l1_q , \sc4_imAck/mxl/muxout , 
        \sc3_wbAck/l1_q , \sc3_wbAck/mxl/muxout , \sc_dm/intI0 , \sc_dm/scn0 , 
        \sc_dm/intI1 , \sc_dm/scn1 , \sc_dm/intI2 , \sc_dm/scn2 , 
        \sc_dm/intI3 , \sc_dm/scn3 , \sc_dm/intI4 , \sc_dm/l4_m/muxout , 
        \sc_dm/l3_m/muxout , \sc_dm/l2_m/muxout , \sc_dm/l1_m/muxout , 
        \sc_dm/l0_m/muxout , \sc_im/intI0 , \sc_im/scn0 , \sc_im/intI1 , 
        \sc_im/scn1 , \sc_im/intI2 , \sc_im/scn2 , \sc_im/intI3 , \sc_im/scn3 , 
        \sc_im/intI4 , \sc_im/l4_m/muxout , \sc_im/l3_m/muxout , 
        \sc_im/l2_m/muxout , \sc_im/l1_m/muxout , \sc_im/l0_m/muxout , 
        \sc_wb/intI0 , \sc_wb/scn0 , \sc_wb/intI1 , \sc_wb/scn1 , 
        \sc_wb/intI2 , \sc_wb/scn2 , \sc_wb/intI3 , \sc_wb/scn3 , 
        \sc_wb/intI4 , \sc_wb/l4_m/muxout , \sc_wb/l3_m/muxout , 
        \sc_wb/l2_m/muxout , \sc_wb/l1_m/muxout , \sc_wb/l0_m/muxout , 
        \sc_dp/scn1 , \sc_dp/scn2 , \sc_dp/scn3 , \sc_dp/scn4 , 
        \sc_dp/sl4/l1_q , \sc_dp/sl4/mxl/muxout , \sc_dp/sl3/l1_q , 
        \sc_dp/sl3/mxl/muxout , \sc_dp/sl2/l1_q , \sc_dp/sl2/mxl/muxout , 
        \sc_dp/sl1/l1_q , \sc_dp/sl1/mxl/muxout , \sc_dp/sl0/l1_q , 
        \sc_dp/sl0/mxl/muxout , \sc_tic/scn1 , \sc_tic/scn2 , \sc_tic/scn3 , 
        \sc_tic/scn4 , \sc_tic/sl4/l1_q , \sc_tic/sl4/mxl/muxout , 
        \sc_tic/sl3/l1_q , \sc_tic/sl3/mxl/muxout , \sc_tic/sl2/l1_q , 
        \sc_tic/sl2/mxl/muxout , \sc_tic/sl1/l1_q , \sc_tic/sl1/mxl/muxout , 
        \sc_tic/sl0/l1_q , \sc_tic/sl0/mxl/muxout , \sc_ip/scn1 , \sc_ip/scn2 , 
        \sc_ip/scn3 , \sc_ip/scn4 , \sc_ip/sl4/l1_q , \sc_ip/sl4/mxl/muxout , 
        \sc_ip/sl3/l1_q , \sc_ip/sl3/mxl/muxout , \sc_ip/sl2/l1_q , 
        \sc_ip/sl2/mxl/muxout , \sc_ip/sl1/l1_q , \sc_ip/sl1/mxl/muxout , 
        \sc_ip/sl0/l1_q , \sc_ip/sl0/mxl/muxout , n1, n2, n3, n4, n5, n6, n7, 
        n8, n9, n10, n11, n12, n13, n14, n15;
    comm_fab fab1 ( .nrst(nrst), .I_port_eop_i(I_port_eop_i_sc), .I_port_d0_i(
        I_port_d0_i_sc), .I_port_d1_i(I_port_d1_i_sc), .I_port_d2_i(
        I_port_d2_i_sc), .I_port_d3_i(I_port_d3_i_sc), .I_port_ack(I_port_ack), 
        .TIC_eop_i(TIC_eop_i_sc), .TIC_d0_i(TIC_d0_i_sc), .TIC_d1_i(
        TIC_d1_i_sc), .TIC_d2_i(TIC_d2_i_sc), .TIC_d3_i(TIC_d3_i_sc), 
        .TIC_ack(TIC_ack), .D_port_eop_i(D_port_eop_i_sc), .D_port_d0_i(
        D_port_d0_i_sc), .D_port_d1_i(D_port_d1_i_sc), .D_port_d2_i(
        D_port_d2_i_sc), .D_port_d3_i(D_port_d3_i_sc), .D_port_ack(D_port_ack), 
        .BC_eop_i(BC_eop_i), .BC_d0_i(BC_d0_i), .BC_d1_i(BC_d1_i), .BC_d2_i(
        BC_d2_i), .BC_d3_i(BC_d3_i), .BC_ack(BC_ack), .WB_eop_i(WB_eop_i), 
        .WB_d0_i(WB_d0_i), .WB_d1_i(WB_d1_i), .WB_d2_i(WB_d2_i), .WB_d3_i(
        WB_d3_i), .WB_ack(WB_ack_sc), .IMEM_eop_i(IMEM_eop_i), .IMEM_d0_i(
        IMEM_d0_i), .IMEM_d1_i(IMEM_d1_i), .IMEM_d2_i(IMEM_d2_i), .IMEM_d3_i(
        IMEM_d3_i), .IMEM_ack(IMEM_ack_sc), .DMEM_eop_i(DMEM_eop_i), 
        .DMEM_d0_i(DMEM_d0_i), .DMEM_d1_i(DMEM_d1_i), .DMEM_d2_i(DMEM_d2_i), 
        .DMEM_d3_i(DMEM_d3_i), .DMEM_ack(DMEM_ack_sc), .test_si(\scan[6] ), 
        .test_so(\scan[7] ), .test_se(n13), .phi1(n9), .phi2(n5), .phi3(n2) );
    latn_1 sc10_s_ipAck ( .q(\scan[11] ), .d(scan_m10), .g(n7) );
    latn_1 sc11_s_ticAck ( .q(\scan[12] ), .d(scan_m11), .g(n4) );
    latn_1 sc12_s_dpAck ( .q(test_so), .d(scan_m12), .g(n6) );
    mux2_1 \sc12_m_dpAck/mux  ( .x(\sc12_m_dpAck/muxout ), .d0(D_port_ack), 
        .sl(n15), .d1(\scan[12] ) );
    latn_1 \sc12_m_dpAck/lph1  ( .q(scan_m12), .d(\sc12_m_dpAck/muxout ), .g(
        n11) );
    mux2_1 \sc11_m_ticAck/mux  ( .x(\sc11_m_ticAck/muxout ), .d0(TIC_ack), 
        .sl(n14), .d1(\scan[11] ) );
    latn_1 \sc11_m_ticAck/lph1  ( .q(scan_m11), .d(\sc11_m_ticAck/muxout ), 
        .g(n8) );
    mux2_1 \sc10_m_ipAck/mux  ( .x(\sc10_m_ipAck/muxout ), .d0(I_port_ack), 
        .sl(n14), .d1(\scan[10] ) );
    latn_1 \sc10_m_ipAck/lph1  ( .q(scan_m10), .d(\sc10_m_ipAck/muxout ), .g(
        n10) );
    latn_1 \sc5_dmAck/lph3  ( .q(DMEM_ack_sc), .d(\sc5_dmAck/l1_q ), .g(n1) );
    latn_1 \sc5_dmAck/lph2  ( .q(\scan[6] ), .d(\sc5_dmAck/l1_q ), .g(n7) );
    mux2_1 \sc5_dmAck/mxl/mux  ( .x(\sc5_dmAck/mxl/muxout ), .d0(DMEM_ack), 
        .sl(n15), .d1(\scan[5] ) );
    latn_1 \sc5_dmAck/mxl/lph1  ( .q(\sc5_dmAck/l1_q ), .d(
        \sc5_dmAck/mxl/muxout ), .g(n10) );
    latn_1 \sc4_imAck/lph3  ( .q(IMEM_ack_sc), .d(\sc4_imAck/l1_q ), .g(n1) );
    latn_1 \sc4_imAck/lph2  ( .q(\scan[5] ), .d(\sc4_imAck/l1_q ), .g(n4) );
    mux2_1 \sc4_imAck/mxl/mux  ( .x(\sc4_imAck/mxl/muxout ), .d0(IMEM_ack), 
        .sl(n12), .d1(\scan[4] ) );
    latn_1 \sc4_imAck/mxl/lph1  ( .q(\sc4_imAck/l1_q ), .d(
        \sc4_imAck/mxl/muxout ), .g(n8) );
    latn_1 \sc3_wbAck/lph3  ( .q(WB_ack_sc), .d(\sc3_wbAck/l1_q ), .g(n1) );
    latn_1 \sc3_wbAck/lph2  ( .q(\scan[4] ), .d(\sc3_wbAck/l1_q ), .g(n6) );
    mux2_1 \sc3_wbAck/mxl/mux  ( .x(\sc3_wbAck/mxl/muxout ), .d0(WB_ack), .sl(
        n12), .d1(\scan[3] ) );
    latn_1 \sc3_wbAck/mxl/lph1  ( .q(\sc3_wbAck/l1_q ), .d(
        \sc3_wbAck/mxl/muxout ), .g(n11) );
    latn_1 \sc_dm/l4_s  ( .q(\scan[10] ), .d(\sc_dm/intI4 ), .g(n7) );
    latn_1 \sc_dm/l3_s  ( .q(\sc_dm/scn3 ), .d(\sc_dm/intI3 ), .g(n4) );
    latn_1 \sc_dm/l2_s  ( .q(\sc_dm/scn2 ), .d(\sc_dm/intI2 ), .g(n6) );
    latn_1 \sc_dm/l1_s  ( .q(\sc_dm/scn1 ), .d(\sc_dm/intI1 ), .g(n7) );
    latn_1 \sc_dm/l0_s  ( .q(\sc_dm/scn0 ), .d(\sc_dm/intI0 ), .g(n4) );
    mux2_1 \sc_dm/l4_m/mux  ( .x(\sc_dm/l4_m/muxout ), .d0(DMEM_d3_i), .sl(n12
        ), .d1(\sc_dm/scn3 ) );
    latn_1 \sc_dm/l4_m/lph1  ( .q(\sc_dm/intI4 ), .d(\sc_dm/l4_m/muxout ), .g(
        n8) );
    mux2_1 \sc_dm/l3_m/mux  ( .x(\sc_dm/l3_m/muxout ), .d0(DMEM_d2_i), .sl(n15
        ), .d1(\sc_dm/scn2 ) );
    latn_1 \sc_dm/l3_m/lph1  ( .q(\sc_dm/intI3 ), .d(\sc_dm/l3_m/muxout ), .g(
        n11) );
    mux2_1 \sc_dm/l2_m/mux  ( .x(\sc_dm/l2_m/muxout ), .d0(DMEM_d1_i), .sl(n14
        ), .d1(\sc_dm/scn1 ) );
    latn_1 \sc_dm/l2_m/lph1  ( .q(\sc_dm/intI2 ), .d(\sc_dm/l2_m/muxout ), .g(
        n10) );
    mux2_1 \sc_dm/l1_m/mux  ( .x(\sc_dm/l1_m/muxout ), .d0(DMEM_d0_i), .sl(n12
        ), .d1(\sc_dm/scn0 ) );
    latn_1 \sc_dm/l1_m/lph1  ( .q(\sc_dm/intI1 ), .d(\sc_dm/l1_m/muxout ), .g(
        n8) );
    mux2_1 \sc_dm/l0_m/mux  ( .x(\sc_dm/l0_m/muxout ), .d0(DMEM_eop_i), .sl(
        n15), .d1(\scan[9] ) );
    latn_1 \sc_dm/l0_m/lph1  ( .q(\sc_dm/intI0 ), .d(\sc_dm/l0_m/muxout ), .g(
        n11) );
    latn_1 \sc_im/l4_s  ( .q(\scan[9] ), .d(\sc_im/intI4 ), .g(n4) );
    latn_1 \sc_im/l3_s  ( .q(\sc_im/scn3 ), .d(\sc_im/intI3 ), .g(n6) );
    latn_1 \sc_im/l2_s  ( .q(\sc_im/scn2 ), .d(\sc_im/intI2 ), .g(n7) );
    latn_1 \sc_im/l1_s  ( .q(\sc_im/scn1 ), .d(\sc_im/intI1 ), .g(n4) );
    latn_1 \sc_im/l0_s  ( .q(\sc_im/scn0 ), .d(\sc_im/intI0 ), .g(n6) );
    mux2_1 \sc_im/l4_m/mux  ( .x(\sc_im/l4_m/muxout ), .d0(IMEM_d3_i), .sl(n14
        ), .d1(\sc_im/scn3 ) );
    latn_1 \sc_im/l4_m/lph1  ( .q(\sc_im/intI4 ), .d(\sc_im/l4_m/muxout ), .g(
        n10) );
    mux2_1 \sc_im/l3_m/mux  ( .x(\sc_im/l3_m/muxout ), .d0(IMEM_d2_i), .sl(n12
        ), .d1(\sc_im/scn2 ) );
    latn_1 \sc_im/l3_m/lph1  ( .q(\sc_im/intI3 ), .d(\sc_im/l3_m/muxout ), .g(
        n8) );
    mux2_1 \sc_im/l2_m/mux  ( .x(\sc_im/l2_m/muxout ), .d0(IMEM_d1_i), .sl(n15
        ), .d1(\sc_im/scn1 ) );
    latn_1 \sc_im/l2_m/lph1  ( .q(\sc_im/intI2 ), .d(\sc_im/l2_m/muxout ), .g(
        n11) );
    mux2_1 \sc_im/l1_m/mux  ( .x(\sc_im/l1_m/muxout ), .d0(IMEM_d0_i), .sl(n14
        ), .d1(\sc_im/scn0 ) );
    latn_1 \sc_im/l1_m/lph1  ( .q(\sc_im/intI1 ), .d(\sc_im/l1_m/muxout ), .g(
        n10) );
    mux2_1 \sc_im/l0_m/mux  ( .x(\sc_im/l0_m/muxout ), .d0(IMEM_eop_i), .sl(
        n12), .d1(\scan[8] ) );
    latn_1 \sc_im/l0_m/lph1  ( .q(\sc_im/intI0 ), .d(\sc_im/l0_m/muxout ), .g(
        n8) );
    latn_1 \sc_wb/l4_s  ( .q(\scan[8] ), .d(\sc_wb/intI4 ), .g(n6) );
    latn_1 \sc_wb/l3_s  ( .q(\sc_wb/scn3 ), .d(\sc_wb/intI3 ), .g(n7) );
    latn_1 \sc_wb/l2_s  ( .q(\sc_wb/scn2 ), .d(\sc_wb/intI2 ), .g(n4) );
    latn_1 \sc_wb/l1_s  ( .q(\sc_wb/scn1 ), .d(\sc_wb/intI1 ), .g(n6) );
    latn_1 \sc_wb/l0_s  ( .q(\sc_wb/scn0 ), .d(\sc_wb/intI0 ), .g(n7) );
    mux2_1 \sc_wb/l4_m/mux  ( .x(\sc_wb/l4_m/muxout ), .d0(WB_d3_i), .sl(n15), 
        .d1(\sc_wb/scn3 ) );
    latn_1 \sc_wb/l4_m/lph1  ( .q(\sc_wb/intI4 ), .d(\sc_wb/l4_m/muxout ), .g(
        n11) );
    mux2_1 \sc_wb/l3_m/mux  ( .x(\sc_wb/l3_m/muxout ), .d0(WB_d2_i), .sl(n15), 
        .d1(\sc_wb/scn2 ) );
    latn_1 \sc_wb/l3_m/lph1  ( .q(\sc_wb/intI3 ), .d(\sc_wb/l3_m/muxout ), .g(
        n10) );
    mux2_1 \sc_wb/l2_m/mux  ( .x(\sc_wb/l2_m/muxout ), .d0(WB_d1_i), .sl(n14), 
        .d1(\sc_wb/scn1 ) );
    latn_1 \sc_wb/l2_m/lph1  ( .q(\sc_wb/intI2 ), .d(\sc_wb/l2_m/muxout ), .g(
        n8) );
    mux2_1 \sc_wb/l1_m/mux  ( .x(\sc_wb/l1_m/muxout ), .d0(WB_d0_i), .sl(n12), 
        .d1(\sc_wb/scn0 ) );
    latn_1 \sc_wb/l1_m/lph1  ( .q(\sc_wb/intI1 ), .d(\sc_wb/l1_m/muxout ), .g(
        n11) );
    mux2_1 \sc_wb/l0_m/mux  ( .x(\sc_wb/l0_m/muxout ), .d0(WB_eop_i), .sl(n15), 
        .d1(\scan[7] ) );
    latn_1 \sc_wb/l0_m/lph1  ( .q(\sc_wb/intI0 ), .d(\sc_wb/l0_m/muxout ), .g(
        n10) );
    latn_1 \sc_dp/sl4/lph3  ( .q(D_port_d3_i_sc), .d(\sc_dp/sl4/l1_q ), .g(n3)
         );
    latn_1 \sc_dp/sl4/lph2  ( .q(\scan[3] ), .d(\sc_dp/sl4/l1_q ), .g(n4) );
    mux2_1 \sc_dp/sl4/mxl/mux  ( .x(\sc_dp/sl4/mxl/muxout ), .d0(D_port_d3_i), 
        .sl(n14), .d1(\sc_dp/scn4 ) );
    latn_1 \sc_dp/sl4/mxl/lph1  ( .q(\sc_dp/sl4/l1_q ), .d(
        \sc_dp/sl4/mxl/muxout ), .g(n8) );
    latn_1 \sc_dp/sl3/lph3  ( .q(D_port_d2_i_sc), .d(\sc_dp/sl3/l1_q ), .g(n3)
         );
    latn_1 \sc_dp/sl3/lph2  ( .q(\sc_dp/scn4 ), .d(\sc_dp/sl3/l1_q ), .g(n7)
         );
    mux2_1 \sc_dp/sl3/mxl/mux  ( .x(\sc_dp/sl3/mxl/muxout ), .d0(D_port_d2_i), 
        .sl(n12), .d1(\sc_dp/scn3 ) );
    latn_1 \sc_dp/sl3/mxl/lph1  ( .q(\sc_dp/sl3/l1_q ), .d(
        \sc_dp/sl3/mxl/muxout ), .g(n11) );
    latn_1 \sc_dp/sl2/lph3  ( .q(D_port_d1_i_sc), .d(\sc_dp/sl2/l1_q ), .g(n3)
         );
    latn_1 \sc_dp/sl2/lph2  ( .q(\sc_dp/scn3 ), .d(\sc_dp/sl2/l1_q ), .g(n6)
         );
    mux2_1 \sc_dp/sl2/mxl/mux  ( .x(\sc_dp/sl2/mxl/muxout ), .d0(D_port_d1_i), 
        .sl(n15), .d1(\sc_dp/scn2 ) );
    latn_1 \sc_dp/sl2/mxl/lph1  ( .q(\sc_dp/sl2/l1_q ), .d(
        \sc_dp/sl2/mxl/muxout ), .g(n10) );
    latn_1 \sc_dp/sl1/lph3  ( .q(D_port_d0_i_sc), .d(\sc_dp/sl1/l1_q ), .g(n3)
         );
    latn_1 \sc_dp/sl1/lph2  ( .q(\sc_dp/scn2 ), .d(\sc_dp/sl1/l1_q ), .g(n7)
         );
    mux2_1 \sc_dp/sl1/mxl/mux  ( .x(\sc_dp/sl1/mxl/muxout ), .d0(D_port_d0_i), 
        .sl(n12), .d1(\sc_dp/scn1 ) );
    latn_1 \sc_dp/sl1/mxl/lph1  ( .q(\sc_dp/sl1/l1_q ), .d(
        \sc_dp/sl1/mxl/muxout ), .g(n11) );
    latn_1 \sc_dp/sl0/lph3  ( .q(D_port_eop_i_sc), .d(\sc_dp/sl0/l1_q ), .g(n3
        ) );
    latn_1 \sc_dp/sl0/lph2  ( .q(\sc_dp/scn1 ), .d(\sc_dp/sl0/l1_q ), .g(n4)
         );
    mux2_1 \sc_dp/sl0/mxl/mux  ( .x(\sc_dp/sl0/mxl/muxout ), .d0(D_port_eop_i), 
        .sl(n12), .d1(\scan[2] ) );
    latn_1 \sc_dp/sl0/mxl/lph1  ( .q(\sc_dp/sl0/l1_q ), .d(
        \sc_dp/sl0/mxl/muxout ), .g(n8) );
    latn_1 \sc_tic/sl4/lph3  ( .q(TIC_d3_i_sc), .d(\sc_tic/sl4/l1_q ), .g(n3)
         );
    latn_1 \sc_tic/sl4/lph2  ( .q(\scan[2] ), .d(\sc_tic/sl4/l1_q ), .g(n6) );
    mux2_1 \sc_tic/sl4/mxl/mux  ( .x(\sc_tic/sl4/mxl/muxout ), .d0(TIC_d3_i), 
        .sl(n14), .d1(\sc_tic/scn4 ) );
    latn_1 \sc_tic/sl4/mxl/lph1  ( .q(\sc_tic/sl4/l1_q ), .d(
        \sc_tic/sl4/mxl/muxout ), .g(n10) );
    latn_1 \sc_tic/sl3/lph3  ( .q(TIC_d2_i_sc), .d(\sc_tic/sl3/l1_q ), .g(n3)
         );
    latn_1 \sc_tic/sl3/lph2  ( .q(\sc_tic/scn4 ), .d(\sc_tic/sl3/l1_q ), .g(n7
        ) );
    mux2_1 \sc_tic/sl3/mxl/mux  ( .x(\sc_tic/sl3/mxl/muxout ), .d0(TIC_d2_i), 
        .sl(n15), .d1(\sc_tic/scn3 ) );
    latn_1 \sc_tic/sl3/mxl/lph1  ( .q(\sc_tic/sl3/l1_q ), .d(
        \sc_tic/sl3/mxl/muxout ), .g(n11) );
    latn_1 \sc_tic/sl2/lph3  ( .q(TIC_d1_i_sc), .d(\sc_tic/sl2/l1_q ), .g(n3)
         );
    latn_1 \sc_tic/sl2/lph2  ( .q(\sc_tic/scn3 ), .d(\sc_tic/sl2/l1_q ), .g(n4
        ) );
    mux2_1 \sc_tic/sl2/mxl/mux  ( .x(\sc_tic/sl2/mxl/muxout ), .d0(TIC_d1_i), 
        .sl(n14), .d1(\sc_tic/scn2 ) );
    latn_1 \sc_tic/sl2/mxl/lph1  ( .q(\sc_tic/sl2/l1_q ), .d(
        \sc_tic/sl2/mxl/muxout ), .g(n8) );
    latn_1 \sc_tic/sl1/lph3  ( .q(TIC_d0_i_sc), .d(\sc_tic/sl1/l1_q ), .g(n3)
         );
    latn_1 \sc_tic/sl1/lph2  ( .q(\sc_tic/scn2 ), .d(\sc_tic/sl1/l1_q ), .g(n7
        ) );
    mux2_1 \sc_tic/sl1/mxl/mux  ( .x(\sc_tic/sl1/mxl/muxout ), .d0(TIC_d0_i), 
        .sl(n15), .d1(\sc_tic/scn1 ) );
    latn_1 \sc_tic/sl1/mxl/lph1  ( .q(\sc_tic/sl1/l1_q ), .d(
        \sc_tic/sl1/mxl/muxout ), .g(n11) );
    latn_1 \sc_tic/sl0/lph3  ( .q(TIC_eop_i_sc), .d(\sc_tic/sl0/l1_q ), .g(n1)
         );
    latn_1 \sc_tic/sl0/lph2  ( .q(\sc_tic/scn1 ), .d(\sc_tic/sl0/l1_q ), .g(n7
        ) );
    mux2_1 \sc_tic/sl0/mxl/mux  ( .x(\sc_tic/sl0/mxl/muxout ), .d0(TIC_eop_i), 
        .sl(n12), .d1(\scan[1] ) );
    latn_1 \sc_tic/sl0/mxl/lph1  ( .q(\sc_tic/sl0/l1_q ), .d(
        \sc_tic/sl0/mxl/muxout ), .g(n11) );
    latn_1 \sc_ip/sl4/lph3  ( .q(I_port_d3_i_sc), .d(\sc_ip/sl4/l1_q ), .g(n1)
         );
    latn_1 \sc_ip/sl4/lph2  ( .q(\scan[1] ), .d(\sc_ip/sl4/l1_q ), .g(n4) );
    mux2_1 \sc_ip/sl4/mxl/mux  ( .x(\sc_ip/sl4/mxl/muxout ), .d0(I_port_d3_i), 
        .sl(n12), .d1(\sc_ip/scn4 ) );
    latn_1 \sc_ip/sl4/mxl/lph1  ( .q(\sc_ip/sl4/l1_q ), .d(
        \sc_ip/sl4/mxl/muxout ), .g(n8) );
    latn_1 \sc_ip/sl3/lph3  ( .q(I_port_d2_i_sc), .d(\sc_ip/sl3/l1_q ), .g(n1)
         );
    latn_1 \sc_ip/sl3/lph2  ( .q(\sc_ip/scn4 ), .d(\sc_ip/sl3/l1_q ), .g(n6)
         );
    mux2_1 \sc_ip/sl3/mxl/mux  ( .x(\sc_ip/sl3/mxl/muxout ), .d0(I_port_d2_i), 
        .sl(n15), .d1(\sc_ip/scn3 ) );
    latn_1 \sc_ip/sl3/mxl/lph1  ( .q(\sc_ip/sl3/l1_q ), .d(
        \sc_ip/sl3/mxl/muxout ), .g(n10) );
    latn_1 \sc_ip/sl2/lph3  ( .q(I_port_d1_i_sc), .d(\sc_ip/sl2/l1_q ), .g(n1)
         );
    latn_1 \sc_ip/sl2/lph2  ( .q(\sc_ip/scn3 ), .d(\sc_ip/sl2/l1_q ), .g(n6)
         );
    mux2_1 \sc_ip/sl2/mxl/mux  ( .x(\sc_ip/sl2/mxl/muxout ), .d0(I_port_d1_i), 
        .sl(n14), .d1(\sc_ip/scn2 ) );
    latn_1 \sc_ip/sl2/mxl/lph1  ( .q(\sc_ip/sl2/l1_q ), .d(
        \sc_ip/sl2/mxl/muxout ), .g(n10) );
    latn_1 \sc_ip/sl1/lph3  ( .q(I_port_d0_i_sc), .d(\sc_ip/sl1/l1_q ), .g(n1)
         );
    latn_1 \sc_ip/sl1/lph2  ( .q(\sc_ip/scn2 ), .d(\sc_ip/sl1/l1_q ), .g(n4)
         );
    mux2_1 \sc_ip/sl1/mxl/mux  ( .x(\sc_ip/sl1/mxl/muxout ), .d0(I_port_d0_i), 
        .sl(n14), .d1(\sc_ip/scn1 ) );
    latn_1 \sc_ip/sl1/mxl/lph1  ( .q(\sc_ip/sl1/l1_q ), .d(
        \sc_ip/sl1/mxl/muxout ), .g(n8) );
    latn_1 \sc_ip/sl0/lph3  ( .q(I_port_eop_i_sc), .d(\sc_ip/sl0/l1_q ), .g(n1
        ) );
    latn_1 \sc_ip/sl0/lph2  ( .q(\sc_ip/scn1 ), .d(\sc_ip/sl0/l1_q ), .g(n6)
         );
    mux2_1 \sc_ip/sl0/mxl/mux  ( .x(\sc_ip/sl0/mxl/muxout ), .d0(I_port_eop_i), 
        .sl(n14), .d1(test_si) );
    latn_1 \sc_ip/sl0/mxl/lph1  ( .q(\sc_ip/sl0/l1_q ), .d(
        \sc_ip/sl0/mxl/muxout ), .g(n10) );
    buf_3 U1 ( .x(n13), .a(test_se) );
    buf_1 U2 ( .x(n1), .a(phi3) );
    buf_1 U3 ( .x(n3), .a(phi3) );
    buf_3 U4 ( .x(n2), .a(phi3) );
    buf_3 U5 ( .x(n4), .a(phi2) );
    buf_3 U6 ( .x(n7), .a(phi2) );
    buf_3 U7 ( .x(n5), .a(phi2) );
    buf_3 U8 ( .x(n6), .a(phi2) );
    buf_3 U9 ( .x(n8), .a(phi1) );
    buf_3 U10 ( .x(n11), .a(phi1) );
    buf_3 U11 ( .x(n9), .a(phi1) );
    buf_3 U12 ( .x(n10), .a(phi1) );
    buf_3 U13 ( .x(n12), .a(test_se) );
    buf_3 U14 ( .x(n15), .a(test_se) );
    buf_3 U15 ( .x(n14), .a(test_se) );
endmodule


module chain_router10 ( eop_i, d0_i, d1_i, d2_i, d3_i, ack_i, eop_ox, d0_ox, 
    d1_ox, d2_ox, d3_ox, ack_ox, eop_oy, d0_oy, d1_oy, d2_oy, d3_oy, ack_oy, 
    nrst, test_si, test_se, test_so, phi1, phi2, phi3 );
input  eop_i, d0_i, d1_i, d2_i, d3_i, ack_ox, ack_oy, nrst, test_si, test_se, 
    phi1, phi2, phi3;
output ack_i, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, eop_oy, d0_oy, d1_oy, d2_oy, 
    d3_oy, test_so;
    wire \scan[2] , \scan[3] , ackx_l, nack_x, sx, acky_l, nack_y, sy, 
        \scan[0] , qa, qa_l, nroutex, routeAckx, nrouteAckx, qx, nqx, neopxy, 
        \scan[1] , sx_pl, nroutey, routeAcky, nrouteAcky, qy, nqy, sy_pl, rst, 
        n10, n11, n12, n1, n2, n3, n4, n5, n6, n7, n8, \cy/__tmp99/nr , 
        \cy/__tmp99/nd , \cx/__tmp99/nr , \cx/__tmp99/nd , \cye/nr , \cye/nd , 
        \cye/n2 , \cy3/__tmp99/loop , \cy2/__tmp99/loop , \cy1/__tmp99/loop , 
        \cy0/__tmp99/loop , \cxe/nr , \cxe/nd , \cxe/n2 , \cx3/__tmp99/loop , 
        \cx2/__tmp99/loop , \cx1/__tmp99/loop , \cx0/__tmp99/loop , 
        \sl_sy/l1_q , \sl_sy/mxl/muxout , \sl_sx/l1_q , \sl_sx/mxl/muxout , 
        \sl_qa/l1_q , \sl_qa/mxl/muxout , \slAcky/l1_q , \slAcky/mxl/muxout , 
        \slAckx/l1_q , \slAckx/mxl/muxout ;
    inv_1 U0 ( .x(rst), .a(nrst) );
    nor2_2 U5 ( .x(nack_x), .a(ackx_l), .b(rst) );
    nor2_2 U4 ( .x(nack_y), .a(acky_l), .b(rst) );
    nand4_1 U1 ( .x(ack_i), .a(n10), .b(n11), .c(n12), .d(neopxy) );
    and4_1 U8 ( .x(n10), .a(n1), .b(n2), .c(n3), .d(n4) );
    inv_1 U10 ( .x(n1), .a(d0_oy) );
    inv_1 U11 ( .x(n2), .a(d1_oy) );
    inv_1 U14 ( .x(n3), .a(d2_oy) );
    inv_1 U16 ( .x(n4), .a(d3_oy) );
    and4_1 U9 ( .x(n11), .a(n5), .b(n6), .c(n7), .d(n8) );
    inv_1 U17 ( .x(n5), .a(d0_ox) );
    inv_1 U18 ( .x(n6), .a(d1_ox) );
    inv_1 U19 ( .x(n7), .a(d2_ox) );
    inv_1 U20 ( .x(n8), .a(d3_ox) );
    nor2_1 U7 ( .x(n12), .a(nrouteAckx), .b(nrouteAcky) );
    nor2_1 U6 ( .x(neopxy), .a(eop_oy), .b(eop_ox) );
    nor2_1 U3 ( .x(nroutex), .a(d3_i), .b(d1_i) );
    nor2_1 U2 ( .x(nroutey), .a(d2_i), .b(d0_i) );
    nand2_1 U12 ( .x(qa), .a(nqx), .b(nqy) );
    nor2i_1 U15 ( .x(sx_pl), .a(qx), .b(nrouteAckx) );
    nor2i_1 U13 ( .x(sy_pl), .a(qy), .b(nrouteAcky) );
    inv_1 \cy/U1  ( .x(nrouteAcky), .a(routeAcky) );
    nor2_1 \cy/__tmp99/U1  ( .x(\cy/__tmp99/nr ), .a(nroutey), .b(qa_l) );
    nand2_1 \cy/__tmp99/U2  ( .x(\cy/__tmp99/nd ), .a(nroutey), .b(qa_l) );
    oai211_1 \cy/__tmp99/U3  ( .x(routeAcky), .a(nrouteAcky), .b(
        \cy/__tmp99/nr ), .c(\cy/__tmp99/nd ), .d(nrst) );
    inv_1 \cx/U1  ( .x(nrouteAckx), .a(routeAckx) );
    nor2_1 \cx/__tmp99/U1  ( .x(\cx/__tmp99/nr ), .a(nroutex), .b(qa_l) );
    nand2_1 \cx/__tmp99/U2  ( .x(\cx/__tmp99/nd ), .a(nroutex), .b(qa_l) );
    oai211_1 \cx/__tmp99/U3  ( .x(routeAckx), .a(nrouteAckx), .b(
        \cx/__tmp99/nr ), .c(\cx/__tmp99/nd ), .d(nrst) );
    nor3_1 \cye/Unr  ( .x(\cye/nr ), .a(eop_i), .b(nack_y), .c(sy) );
    nand3_1 \cye/Und  ( .x(\cye/nd ), .a(eop_i), .b(nack_y), .c(sy) );
    oa21_1 \cye/U1  ( .x(\cye/n2 ), .a(\cye/n2 ), .b(\cye/nr ), .c(\cye/nd )
         );
    inv_1 \cye/U3  ( .x(eop_oy), .a(\cye/n2 ) );
    ao31_1 \cy3/__tmp99/aoi  ( .x(\cy3/__tmp99/loop ), .a(d3_i), .b(nack_y), 
        .c(sy), .d(d3_oy) );
    ao31_1 \cy2/__tmp99/aoi  ( .x(\cy2/__tmp99/loop ), .a(d2_i), .b(nack_y), 
        .c(sy), .d(d2_oy) );
    ao31_1 \cy1/__tmp99/aoi  ( .x(\cy1/__tmp99/loop ), .a(d1_i), .b(nack_y), 
        .c(sy), .d(d1_oy) );
    ao31_1 \cy0/__tmp99/aoi  ( .x(\cy0/__tmp99/loop ), .a(d0_i), .b(nack_y), 
        .c(sy), .d(d0_oy) );
    nor3_1 \cxe/Unr  ( .x(\cxe/nr ), .a(eop_i), .b(nack_x), .c(sx) );
    nand3_1 \cxe/Und  ( .x(\cxe/nd ), .a(eop_i), .b(nack_x), .c(sx) );
    oa21_1 \cxe/U1  ( .x(\cxe/n2 ), .a(\cxe/n2 ), .b(\cxe/nr ), .c(\cxe/nd )
         );
    inv_1 \cxe/U3  ( .x(eop_ox), .a(\cxe/n2 ) );
    ao31_1 \cx3/__tmp99/aoi  ( .x(\cx3/__tmp99/loop ), .a(d3_i), .b(nack_x), 
        .c(sx), .d(d3_ox) );
    oa21_1 \cx3/__tmp99/outGate  ( .x(d3_ox), .a(d3_i), .b(nack_x), .c(
        \cx3/__tmp99/loop ) );
    ao31_1 \cx2/__tmp99/aoi  ( .x(\cx2/__tmp99/loop ), .a(d2_i), .b(nack_x), 
        .c(sx), .d(d2_ox) );
    oa21_1 \cx2/__tmp99/outGate  ( .x(d2_ox), .a(d2_i), .b(nack_x), .c(
        \cx2/__tmp99/loop ) );
    ao31_1 \cx1/__tmp99/aoi  ( .x(\cx1/__tmp99/loop ), .a(d1_i), .b(nack_x), 
        .c(sx), .d(d1_ox) );
    oa21_1 \cx1/__tmp99/outGate  ( .x(d1_ox), .a(d1_i), .b(nack_x), .c(
        \cx1/__tmp99/loop ) );
    ao31_1 \cx0/__tmp99/aoi  ( .x(\cx0/__tmp99/loop ), .a(d0_i), .b(nack_x), 
        .c(sx), .d(d0_ox) );
    oa21_1 \cx0/__tmp99/outGate  ( .x(d0_ox), .a(d0_i), .b(nack_x), .c(
        \cx0/__tmp99/loop ) );
    nand3_1 \sry/i0  ( .x(nqy), .a(neopxy), .b(nrst), .c(qy) );
    nand2_1 \sry/i1  ( .x(qy), .a(routeAcky), .b(nqy) );
    nand3_1 \srx/i0  ( .x(nqx), .a(neopxy), .b(nrst), .c(qx) );
    nand2_1 \srx/i1  ( .x(qx), .a(routeAckx), .b(nqx) );
    latn_1 \sl_sy/lph3  ( .q(sy), .d(\sl_sy/l1_q ), .g(phi3) );
    latn_1 \sl_sy/lph2  ( .q(\scan[2] ), .d(\sl_sy/l1_q ), .g(phi2) );
    mux2_1 \sl_sy/mxl/mux  ( .x(\sl_sy/mxl/muxout ), .d0(sy_pl), .sl(test_se), 
        .d1(\scan[1] ) );
    latn_1 \sl_sy/mxl/lph1  ( .q(\sl_sy/l1_q ), .d(\sl_sy/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_sx/lph3  ( .q(sx), .d(\sl_sx/l1_q ), .g(phi3) );
    latn_1 \sl_sx/lph2  ( .q(\scan[1] ), .d(\sl_sx/l1_q ), .g(phi2) );
    mux2_1 \sl_sx/mxl/mux  ( .x(\sl_sx/mxl/muxout ), .d0(sx_pl), .sl(test_se), 
        .d1(\scan[0] ) );
    latn_1 \sl_sx/mxl/lph1  ( .q(\sl_sx/l1_q ), .d(\sl_sx/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_qa/lph3  ( .q(qa_l), .d(\sl_qa/l1_q ), .g(phi3) );
    latn_1 \sl_qa/lph2  ( .q(\scan[0] ), .d(\sl_qa/l1_q ), .g(phi2) );
    mux2_1 \sl_qa/mxl/mux  ( .x(\sl_qa/mxl/muxout ), .d0(qa), .sl(test_se), 
        .d1(test_si) );
    latn_1 \sl_qa/mxl/lph1  ( .q(\sl_qa/l1_q ), .d(\sl_qa/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAcky/lph3  ( .q(acky_l), .d(\slAcky/l1_q ), .g(phi3) );
    latn_1 \slAcky/lph2  ( .q(test_so), .d(\slAcky/l1_q ), .g(phi2) );
    mux2_1 \slAcky/mxl/mux  ( .x(\slAcky/mxl/muxout ), .d0(ack_oy), .sl(
        test_se), .d1(\scan[3] ) );
    latn_1 \slAcky/mxl/lph1  ( .q(\slAcky/l1_q ), .d(\slAcky/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAckx/lph3  ( .q(ackx_l), .d(\slAckx/l1_q ), .g(phi3) );
    latn_1 \slAckx/lph2  ( .q(\scan[3] ), .d(\slAckx/l1_q ), .g(phi2) );
    mux2_1 \slAckx/mxl/mux  ( .x(\slAckx/mxl/muxout ), .d0(ack_ox), .sl(
        test_se), .d1(\scan[2] ) );
    latn_1 \slAckx/mxl/lph1  ( .q(\slAckx/l1_q ), .d(\slAckx/mxl/muxout ), .g(
        phi1) );
    oa21_2 U21 ( .x(d1_oy), .a(d1_i), .b(nack_y), .c(\cy1/__tmp99/loop ) );
    oa21_2 U22 ( .x(d2_oy), .a(d2_i), .b(nack_y), .c(\cy2/__tmp99/loop ) );
    oa21_2 U23 ( .x(d0_oy), .a(d0_i), .b(nack_y), .c(\cy0/__tmp99/loop ) );
    oa21_2 U24 ( .x(d3_oy), .a(d3_i), .b(nack_y), .c(\cy3/__tmp99/loop ) );
endmodule


module chain_router11 ( eop_i, d0_i, d1_i, d2_i, d3_i, ack_i, eop_ox, d0_ox, 
    d1_ox, d2_ox, d3_ox, ack_ox, eop_oy, d0_oy, d1_oy, d2_oy, d3_oy, ack_oy, 
    nrst, test_si, test_se, test_so, phi1, phi2, phi3 );
input  eop_i, d0_i, d1_i, d2_i, d3_i, ack_ox, ack_oy, nrst, test_si, test_se, 
    phi1, phi2, phi3;
output ack_i, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, eop_oy, d0_oy, d1_oy, d2_oy, 
    d3_oy, test_so;
    wire \scan[2] , \scan[3] , ackx_l, nack_x, sx, acky_l, nack_y, sy, 
        \scan[0] , qa, qa_l, nroutex, routeAckx, nrouteAckx, qx, nqx, neopxy, 
        \scan[1] , sx_pl, nroutey, routeAcky, nrouteAcky, qy, nqy, sy_pl, rst, 
        n10, n11, n12, n1, n2, n3, n4, n5, n6, n7, n8, \cy/__tmp99/nr , 
        \cy/__tmp99/nd , \cx/__tmp99/nr , \cx/__tmp99/nd , \cye/nr , \cye/nd , 
        \cye/n2 , \cy3/__tmp99/loop , \cy2/__tmp99/loop , \cy1/__tmp99/loop , 
        \cy0/__tmp99/loop , \cxe/nr , \cxe/nd , \cxe/n2 , \cx3/__tmp99/loop , 
        \cx2/__tmp99/loop , \cx1/__tmp99/loop , \cx0/__tmp99/loop , 
        \sl_sy/l1_q , \sl_sy/mxl/muxout , \sl_sx/l1_q , \sl_sx/mxl/muxout , 
        \sl_qa/l1_q , \sl_qa/mxl/muxout , \slAcky/l1_q , \slAcky/mxl/muxout , 
        \slAckx/l1_q , \slAckx/mxl/muxout ;
    inv_1 U0 ( .x(rst), .a(nrst) );
    nor2_2 U5 ( .x(nack_x), .a(ackx_l), .b(rst) );
    nor2_2 U4 ( .x(nack_y), .a(acky_l), .b(rst) );
    nand4_1 U1 ( .x(ack_i), .a(n10), .b(n11), .c(n12), .d(neopxy) );
    and4_1 U8 ( .x(n10), .a(n1), .b(n2), .c(n3), .d(n4) );
    inv_1 U10 ( .x(n1), .a(d0_oy) );
    inv_1 U11 ( .x(n2), .a(d1_oy) );
    inv_1 U14 ( .x(n3), .a(d2_oy) );
    inv_1 U16 ( .x(n4), .a(d3_oy) );
    and4_1 U9 ( .x(n11), .a(n5), .b(n6), .c(n7), .d(n8) );
    inv_1 U17 ( .x(n5), .a(d0_ox) );
    inv_1 U18 ( .x(n6), .a(d1_ox) );
    inv_1 U19 ( .x(n7), .a(d2_ox) );
    inv_1 U20 ( .x(n8), .a(d3_ox) );
    nor2_1 U7 ( .x(n12), .a(nrouteAckx), .b(nrouteAcky) );
    nor2_1 U6 ( .x(neopxy), .a(eop_oy), .b(eop_ox) );
    nor2_1 U3 ( .x(nroutex), .a(d3_i), .b(d1_i) );
    nor2_1 U2 ( .x(nroutey), .a(d2_i), .b(d0_i) );
    nand2_1 U12 ( .x(qa), .a(nqx), .b(nqy) );
    nor2i_1 U15 ( .x(sx_pl), .a(qx), .b(nrouteAckx) );
    nor2i_1 U13 ( .x(sy_pl), .a(qy), .b(nrouteAcky) );
    inv_1 \cy/U1  ( .x(nrouteAcky), .a(routeAcky) );
    nor2_1 \cy/__tmp99/U1  ( .x(\cy/__tmp99/nr ), .a(nroutey), .b(qa_l) );
    nand2_1 \cy/__tmp99/U2  ( .x(\cy/__tmp99/nd ), .a(nroutey), .b(qa_l) );
    oai211_1 \cy/__tmp99/U3  ( .x(routeAcky), .a(nrouteAcky), .b(
        \cy/__tmp99/nr ), .c(\cy/__tmp99/nd ), .d(nrst) );
    inv_1 \cx/U1  ( .x(nrouteAckx), .a(routeAckx) );
    nor2_1 \cx/__tmp99/U1  ( .x(\cx/__tmp99/nr ), .a(nroutex), .b(qa_l) );
    nand2_1 \cx/__tmp99/U2  ( .x(\cx/__tmp99/nd ), .a(nroutex), .b(qa_l) );
    oai211_1 \cx/__tmp99/U3  ( .x(routeAckx), .a(nrouteAckx), .b(
        \cx/__tmp99/nr ), .c(\cx/__tmp99/nd ), .d(nrst) );
    nor3_1 \cye/Unr  ( .x(\cye/nr ), .a(eop_i), .b(nack_y), .c(sy) );
    nand3_1 \cye/Und  ( .x(\cye/nd ), .a(eop_i), .b(nack_y), .c(sy) );
    oa21_1 \cye/U1  ( .x(\cye/n2 ), .a(\cye/n2 ), .b(\cye/nr ), .c(\cye/nd )
         );
    inv_1 \cye/U3  ( .x(eop_oy), .a(\cye/n2 ) );
    ao31_1 \cy3/__tmp99/aoi  ( .x(\cy3/__tmp99/loop ), .a(d3_i), .b(nack_y), 
        .c(sy), .d(d3_oy) );
    ao31_1 \cy2/__tmp99/aoi  ( .x(\cy2/__tmp99/loop ), .a(d2_i), .b(nack_y), 
        .c(sy), .d(d2_oy) );
    ao31_1 \cy1/__tmp99/aoi  ( .x(\cy1/__tmp99/loop ), .a(d1_i), .b(nack_y), 
        .c(sy), .d(d1_oy) );
    ao31_1 \cy0/__tmp99/aoi  ( .x(\cy0/__tmp99/loop ), .a(d0_i), .b(nack_y), 
        .c(sy), .d(d0_oy) );
    nor3_1 \cxe/Unr  ( .x(\cxe/nr ), .a(eop_i), .b(nack_x), .c(sx) );
    nand3_1 \cxe/Und  ( .x(\cxe/nd ), .a(eop_i), .b(nack_x), .c(sx) );
    oa21_1 \cxe/U1  ( .x(\cxe/n2 ), .a(\cxe/n2 ), .b(\cxe/nr ), .c(\cxe/nd )
         );
    inv_1 \cxe/U3  ( .x(eop_ox), .a(\cxe/n2 ) );
    ao31_1 \cx3/__tmp99/aoi  ( .x(\cx3/__tmp99/loop ), .a(d3_i), .b(nack_x), 
        .c(sx), .d(d3_ox) );
    ao31_1 \cx2/__tmp99/aoi  ( .x(\cx2/__tmp99/loop ), .a(d2_i), .b(nack_x), 
        .c(sx), .d(d2_ox) );
    ao31_1 \cx1/__tmp99/aoi  ( .x(\cx1/__tmp99/loop ), .a(d1_i), .b(nack_x), 
        .c(sx), .d(d1_ox) );
    ao31_1 \cx0/__tmp99/aoi  ( .x(\cx0/__tmp99/loop ), .a(d0_i), .b(nack_x), 
        .c(sx), .d(d0_ox) );
    nand3_1 \sry/i0  ( .x(nqy), .a(neopxy), .b(nrst), .c(qy) );
    nand2_1 \sry/i1  ( .x(qy), .a(routeAcky), .b(nqy) );
    nand3_1 \srx/i0  ( .x(nqx), .a(neopxy), .b(nrst), .c(qx) );
    nand2_1 \srx/i1  ( .x(qx), .a(routeAckx), .b(nqx) );
    latn_1 \sl_sy/lph3  ( .q(sy), .d(\sl_sy/l1_q ), .g(phi3) );
    latn_1 \sl_sy/lph2  ( .q(\scan[2] ), .d(\sl_sy/l1_q ), .g(phi2) );
    mux2_1 \sl_sy/mxl/mux  ( .x(\sl_sy/mxl/muxout ), .d0(sy_pl), .sl(test_se), 
        .d1(\scan[1] ) );
    latn_1 \sl_sy/mxl/lph1  ( .q(\sl_sy/l1_q ), .d(\sl_sy/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_sx/lph3  ( .q(sx), .d(\sl_sx/l1_q ), .g(phi3) );
    latn_1 \sl_sx/lph2  ( .q(\scan[1] ), .d(\sl_sx/l1_q ), .g(phi2) );
    mux2_1 \sl_sx/mxl/mux  ( .x(\sl_sx/mxl/muxout ), .d0(sx_pl), .sl(test_se), 
        .d1(\scan[0] ) );
    latn_1 \sl_sx/mxl/lph1  ( .q(\sl_sx/l1_q ), .d(\sl_sx/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_qa/lph3  ( .q(qa_l), .d(\sl_qa/l1_q ), .g(phi3) );
    latn_1 \sl_qa/lph2  ( .q(\scan[0] ), .d(\sl_qa/l1_q ), .g(phi2) );
    mux2_1 \sl_qa/mxl/mux  ( .x(\sl_qa/mxl/muxout ), .d0(qa), .sl(test_se), 
        .d1(test_si) );
    latn_1 \sl_qa/mxl/lph1  ( .q(\sl_qa/l1_q ), .d(\sl_qa/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAcky/lph3  ( .q(acky_l), .d(\slAcky/l1_q ), .g(phi3) );
    latn_1 \slAcky/lph2  ( .q(test_so), .d(\slAcky/l1_q ), .g(phi2) );
    mux2_1 \slAcky/mxl/mux  ( .x(\slAcky/mxl/muxout ), .d0(ack_oy), .sl(
        test_se), .d1(\scan[3] ) );
    latn_1 \slAcky/mxl/lph1  ( .q(\slAcky/l1_q ), .d(\slAcky/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAckx/lph3  ( .q(ackx_l), .d(\slAckx/l1_q ), .g(phi3) );
    latn_1 \slAckx/lph2  ( .q(\scan[3] ), .d(\slAckx/l1_q ), .g(phi2) );
    mux2_1 \slAckx/mxl/mux  ( .x(\slAckx/mxl/muxout ), .d0(ack_ox), .sl(
        test_se), .d1(\scan[2] ) );
    latn_1 \slAckx/mxl/lph1  ( .q(\slAckx/l1_q ), .d(\slAckx/mxl/muxout ), .g(
        phi1) );
    oa21_2 U21 ( .x(d3_oy), .a(d3_i), .b(nack_y), .c(\cy3/__tmp99/loop ) );
    oa21_2 U22 ( .x(d2_oy), .a(d2_i), .b(nack_y), .c(\cy2/__tmp99/loop ) );
    oa21_2 U23 ( .x(d1_oy), .a(d1_i), .b(nack_y), .c(\cy1/__tmp99/loop ) );
    oa21_2 U24 ( .x(d0_ox), .a(d0_i), .b(nack_x), .c(\cx0/__tmp99/loop ) );
    oa21_2 U25 ( .x(d2_ox), .a(d2_i), .b(nack_x), .c(\cx2/__tmp99/loop ) );
    oa21_2 U26 ( .x(d3_ox), .a(d3_i), .b(nack_x), .c(\cx3/__tmp99/loop ) );
    oa21_2 U27 ( .x(d1_ox), .a(d1_i), .b(nack_x), .c(\cx1/__tmp99/loop ) );
    oa21_2 U28 ( .x(d0_oy), .a(d0_i), .b(nack_y), .c(\cy0/__tmp99/loop ) );
endmodule


module chain_arbiter10 ( eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, ack_ix, eop_iy, 
    d0_iy, d1_iy, d2_iy, d3_iy, ack_iy, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, 
    eop_oy, d0_oy, d1_oy, d2_oy, d3_oy, ack_oxy, rst, test_si, test_se, 
    test_so, phi1, phi2, phi3 );
input  eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, eop_iy, d0_iy, d1_iy, d2_iy, d3_iy, 
    ack_oxy, rst, test_si, test_se, phi1, phi2, phi3;
output ack_ix, ack_iy, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, eop_oy, d0_oy, 
    d1_oy, d2_oy, d3_oy, test_so;
    wire \scan[1] , \scan[2] , ackx_l, nack_x, sx, acky_l, nack_y, sy, mrx, 
        req_x, mry, req_y, gx, gy, \scan[0] , sx_pl, sy_pl, n1x, n2x, n1y, n2y, 
        n5x, n6x, n5y, n6y, \cye/nr , \cye/nd , \cye/n2 , \cy3/__tmp99/loop , 
        \cy2/__tmp99/loop , \cy1/__tmp99/loop , \cy0/__tmp99/loop , \cxe/nr , 
        \cxe/nd , \cxe/n2 , \cx3/__tmp99/loop , \cx2/__tmp99/loop , 
        \cx1/__tmp99/loop , \cx0/__tmp99/loop , \mtx/gr2 , \mtx/gr1 , \sry/qz , 
        \srx/qz , \sl_sy/l1_q , \sl_sy/mxl/muxout , \sl_sx/l1_q , 
        \sl_sx/mxl/muxout , \slAcky/l1_q , \slAcky/mxl/muxout , \slAckx/l1_q , 
        \slAckx/mxl/muxout ;
    nor2_2 U12 ( .x(nack_x), .a(ackx_l), .b(rst) );
    nand2_1 U4 ( .x(ack_ix), .a(n1x), .b(n2x) );
    nor3_1 U17 ( .x(n1x), .a(d2_ox), .b(d3_ox), .c(d1_ox) );
    nor2_1 U18 ( .x(n2x), .a(eop_ox), .b(d0_ox) );
    nor2_2 U11 ( .x(nack_y), .a(acky_l), .b(rst) );
    nand2_1 U3 ( .x(ack_iy), .a(n1y), .b(n2y) );
    nor3_1 U16 ( .x(n1y), .a(d2_oy), .b(d3_oy), .c(d1_oy) );
    nor2_1 U19 ( .x(n2y), .a(eop_oy), .b(d0_oy) );
    nand2_1 U15 ( .x(req_x), .a(n5x), .b(n6x) );
    nor3_1 U10 ( .x(n5x), .a(d2_ix), .b(d3_ix), .c(d1_ix) );
    nor2_1 U13 ( .x(n6x), .a(eop_ix), .b(d0_ix) );
    nand2_1 U14 ( .x(req_y), .a(n5y), .b(n6y) );
    nor3_1 U9 ( .x(n5y), .a(d2_iy), .b(d3_iy), .c(d1_iy) );
    nor2_1 U20 ( .x(n6y), .a(eop_iy), .b(d0_iy) );
    nor2i_1 U6 ( .x(sx_pl), .a(gx), .b(eop_oy) );
    nor2i_1 U5 ( .x(sy_pl), .a(gy), .b(eop_ox) );
    nor3_1 \cye/Unr  ( .x(\cye/nr ), .a(eop_iy), .b(nack_y), .c(sy) );
    nand3_1 \cye/Und  ( .x(\cye/nd ), .a(eop_iy), .b(nack_y), .c(sy) );
    oa21_1 \cye/U1  ( .x(\cye/n2 ), .a(\cye/n2 ), .b(\cye/nr ), .c(\cye/nd )
         );
    inv_1 \cye/U3  ( .x(eop_oy), .a(\cye/n2 ) );
    ao31_1 \cy3/__tmp99/aoi  ( .x(\cy3/__tmp99/loop ), .a(d3_iy), .b(nack_y), 
        .c(sy), .d(d3_oy) );
    oa21_1 \cy3/__tmp99/outGate  ( .x(d3_oy), .a(d3_iy), .b(nack_y), .c(
        \cy3/__tmp99/loop ) );
    ao31_1 \cy2/__tmp99/aoi  ( .x(\cy2/__tmp99/loop ), .a(d2_iy), .b(nack_y), 
        .c(sy), .d(d2_oy) );
    oa21_1 \cy2/__tmp99/outGate  ( .x(d2_oy), .a(d2_iy), .b(nack_y), .c(
        \cy2/__tmp99/loop ) );
    ao31_1 \cy1/__tmp99/aoi  ( .x(\cy1/__tmp99/loop ), .a(d1_iy), .b(nack_y), 
        .c(sy), .d(d1_oy) );
    oa21_1 \cy1/__tmp99/outGate  ( .x(d1_oy), .a(d1_iy), .b(nack_y), .c(
        \cy1/__tmp99/loop ) );
    ao31_1 \cy0/__tmp99/aoi  ( .x(\cy0/__tmp99/loop ), .a(d0_iy), .b(nack_y), 
        .c(sy), .d(d0_oy) );
    oa21_1 \cy0/__tmp99/outGate  ( .x(d0_oy), .a(d0_iy), .b(nack_y), .c(
        \cy0/__tmp99/loop ) );
    nor3_1 \cxe/Unr  ( .x(\cxe/nr ), .a(eop_ix), .b(nack_x), .c(sx) );
    nand3_1 \cxe/Und  ( .x(\cxe/nd ), .a(eop_ix), .b(nack_x), .c(sx) );
    oa21_1 \cxe/U1  ( .x(\cxe/n2 ), .a(\cxe/n2 ), .b(\cxe/nr ), .c(\cxe/nd )
         );
    inv_1 \cxe/U3  ( .x(eop_ox), .a(\cxe/n2 ) );
    ao31_1 \cx3/__tmp99/aoi  ( .x(\cx3/__tmp99/loop ), .a(d3_ix), .b(nack_x), 
        .c(sx), .d(d3_ox) );
    oa21_1 \cx3/__tmp99/outGate  ( .x(d3_ox), .a(d3_ix), .b(nack_x), .c(
        \cx3/__tmp99/loop ) );
    ao31_1 \cx2/__tmp99/aoi  ( .x(\cx2/__tmp99/loop ), .a(d2_ix), .b(nack_x), 
        .c(sx), .d(d2_ox) );
    oa21_1 \cx2/__tmp99/outGate  ( .x(d2_ox), .a(d2_ix), .b(nack_x), .c(
        \cx2/__tmp99/loop ) );
    ao31_1 \cx1/__tmp99/aoi  ( .x(\cx1/__tmp99/loop ), .a(d1_ix), .b(nack_x), 
        .c(sx), .d(d1_ox) );
    oa21_1 \cx1/__tmp99/outGate  ( .x(d1_ox), .a(d1_ix), .b(nack_x), .c(
        \cx1/__tmp99/loop ) );
    ao31_1 \cx0/__tmp99/aoi  ( .x(\cx0/__tmp99/loop ), .a(d0_ix), .b(nack_x), 
        .c(sx), .d(d0_ox) );
    oa21_1 \cx0/__tmp99/outGate  ( .x(d0_ox), .a(d0_ix), .b(nack_x), .c(
        \cx0/__tmp99/loop ) );
    nand2_1 \mtx/mg2  ( .x(\mtx/gr2 ), .a(mry), .b(\mtx/gr1 ) );
    nand2_1 \mtx/U1  ( .x(\mtx/gr1 ), .a(mrx), .b(\mtx/gr2 ) );
    nor3_1 \mtx/U2  ( .x(gy), .a(\mtx/gr2 ), .b(\mtx/gr2 ), .c(\mtx/gr2 ) );
    nor3_1 \mtx/U3  ( .x(gx), .a(\mtx/gr1 ), .b(\mtx/gr1 ), .c(\mtx/gr1 ) );
    nor2_1 \sry/i1  ( .x(\sry/qz ), .a(req_y), .b(mry) );
    nor2_1 \srx/i1  ( .x(\srx/qz ), .a(req_x), .b(mrx) );
    latn_1 \sl_sy/lph3  ( .q(sy), .d(\sl_sy/l1_q ), .g(phi3) );
    latn_1 \sl_sy/lph2  ( .q(\scan[1] ), .d(\sl_sy/l1_q ), .g(phi2) );
    mux2_1 \sl_sy/mxl/mux  ( .x(\sl_sy/mxl/muxout ), .d0(sy_pl), .sl(test_se), 
        .d1(\scan[0] ) );
    latn_1 \sl_sy/mxl/lph1  ( .q(\sl_sy/l1_q ), .d(\sl_sy/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_sx/lph3  ( .q(sx), .d(\sl_sx/l1_q ), .g(phi3) );
    latn_1 \sl_sx/lph2  ( .q(\scan[0] ), .d(\sl_sx/l1_q ), .g(phi2) );
    mux2_1 \sl_sx/mxl/mux  ( .x(\sl_sx/mxl/muxout ), .d0(sx_pl), .sl(test_se), 
        .d1(test_si) );
    latn_1 \sl_sx/mxl/lph1  ( .q(\sl_sx/l1_q ), .d(\sl_sx/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAcky/lph3  ( .q(acky_l), .d(\slAcky/l1_q ), .g(phi3) );
    latn_1 \slAcky/lph2  ( .q(test_so), .d(\slAcky/l1_q ), .g(phi2) );
    mux2_1 \slAcky/mxl/mux  ( .x(\slAcky/mxl/muxout ), .d0(ack_oxy), .sl(
        test_se), .d1(\scan[2] ) );
    latn_1 \slAcky/mxl/lph1  ( .q(\slAcky/l1_q ), .d(\slAcky/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAckx/lph3  ( .q(ackx_l), .d(\slAckx/l1_q ), .g(phi3) );
    latn_1 \slAckx/lph2  ( .q(\scan[2] ), .d(\slAckx/l1_q ), .g(phi2) );
    mux2_1 \slAckx/mxl/mux  ( .x(\slAckx/mxl/muxout ), .d0(ack_oxy), .sl(
        test_se), .d1(\scan[1] ) );
    latn_1 \slAckx/mxl/lph1  ( .q(\slAckx/l1_q ), .d(\slAckx/mxl/muxout ), .g(
        phi1) );
    nor3_1 U1 ( .x(mry), .a(eop_oy), .b(rst), .c(\sry/qz ) );
    nor3_1 U2 ( .x(mrx), .a(eop_ox), .b(rst), .c(\srx/qz ) );
endmodule


module chain_arbiter11 ( eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, ack_ix, eop_iy, 
    d0_iy, d1_iy, d2_iy, d3_iy, ack_iy, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, 
    eop_oy, d0_oy, d1_oy, d2_oy, d3_oy, ack_oxy, rst, test_si, test_se, 
    test_so, phi1, phi2, phi3 );
input  eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, eop_iy, d0_iy, d1_iy, d2_iy, d3_iy, 
    ack_oxy, rst, test_si, test_se, phi1, phi2, phi3;
output ack_ix, ack_iy, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, eop_oy, d0_oy, 
    d1_oy, d2_oy, d3_oy, test_so;
    wire \scan[1] , \scan[2] , ackx_l, nack_x, sx, acky_l, nack_y, sy, mrx, 
        req_x, mry, req_y, gx, gy, \scan[0] , sx_pl, sy_pl, n1x, n2x, n1y, n2y, 
        n5x, n6x, n5y, n6y, \cye/nr , \cye/nd , \cye/n2 , \cy3/__tmp99/loop , 
        \cy2/__tmp99/loop , \cy1/__tmp99/loop , \cy0/__tmp99/loop , \cxe/nr , 
        \cxe/nd , \cxe/n2 , \cx3/__tmp99/loop , \cx2/__tmp99/loop , 
        \cx1/__tmp99/loop , \cx0/__tmp99/loop , \mtx/gr2 , \mtx/gr1 , \sry/qz , 
        \srx/qz , \sl_sy/l1_q , \sl_sy/mxl/muxout , \sl_sx/l1_q , 
        \sl_sx/mxl/muxout , \slAcky/l1_q , \slAcky/mxl/muxout , \slAckx/l1_q , 
        \slAckx/mxl/muxout ;
    nor2_2 U12 ( .x(nack_x), .a(ackx_l), .b(rst) );
    nand2_1 U4 ( .x(ack_ix), .a(n1x), .b(n2x) );
    nor3_1 U17 ( .x(n1x), .a(d2_ox), .b(d3_ox), .c(d1_ox) );
    nor2_1 U18 ( .x(n2x), .a(eop_ox), .b(d0_ox) );
    nor2_2 U11 ( .x(nack_y), .a(acky_l), .b(rst) );
    nand2_1 U3 ( .x(ack_iy), .a(n1y), .b(n2y) );
    nor3_1 U16 ( .x(n1y), .a(d2_oy), .b(d3_oy), .c(d1_oy) );
    nor2_1 U19 ( .x(n2y), .a(eop_oy), .b(d0_oy) );
    nand2_1 U15 ( .x(req_x), .a(n5x), .b(n6x) );
    nor3_1 U10 ( .x(n5x), .a(d2_ix), .b(d3_ix), .c(d1_ix) );
    nor2_1 U13 ( .x(n6x), .a(eop_ix), .b(d0_ix) );
    nand2_1 U14 ( .x(req_y), .a(n5y), .b(n6y) );
    nor3_1 U9 ( .x(n5y), .a(d2_iy), .b(d3_iy), .c(d1_iy) );
    nor2_1 U20 ( .x(n6y), .a(eop_iy), .b(d0_iy) );
    nor2i_1 U6 ( .x(sx_pl), .a(gx), .b(eop_oy) );
    nor2i_1 U5 ( .x(sy_pl), .a(gy), .b(eop_ox) );
    nor3_1 \cye/Unr  ( .x(\cye/nr ), .a(eop_iy), .b(nack_y), .c(sy) );
    nand3_1 \cye/Und  ( .x(\cye/nd ), .a(eop_iy), .b(nack_y), .c(sy) );
    oa21_1 \cye/U1  ( .x(\cye/n2 ), .a(\cye/n2 ), .b(\cye/nr ), .c(\cye/nd )
         );
    inv_1 \cye/U3  ( .x(eop_oy), .a(\cye/n2 ) );
    ao31_1 \cy3/__tmp99/aoi  ( .x(\cy3/__tmp99/loop ), .a(d3_iy), .b(nack_y), 
        .c(sy), .d(d3_oy) );
    oa21_1 \cy3/__tmp99/outGate  ( .x(d3_oy), .a(d3_iy), .b(nack_y), .c(
        \cy3/__tmp99/loop ) );
    ao31_1 \cy2/__tmp99/aoi  ( .x(\cy2/__tmp99/loop ), .a(d2_iy), .b(nack_y), 
        .c(sy), .d(d2_oy) );
    oa21_1 \cy2/__tmp99/outGate  ( .x(d2_oy), .a(d2_iy), .b(nack_y), .c(
        \cy2/__tmp99/loop ) );
    ao31_1 \cy1/__tmp99/aoi  ( .x(\cy1/__tmp99/loop ), .a(d1_iy), .b(nack_y), 
        .c(sy), .d(d1_oy) );
    oa21_1 \cy1/__tmp99/outGate  ( .x(d1_oy), .a(d1_iy), .b(nack_y), .c(
        \cy1/__tmp99/loop ) );
    ao31_1 \cy0/__tmp99/aoi  ( .x(\cy0/__tmp99/loop ), .a(d0_iy), .b(nack_y), 
        .c(sy), .d(d0_oy) );
    oa21_1 \cy0/__tmp99/outGate  ( .x(d0_oy), .a(d0_iy), .b(nack_y), .c(
        \cy0/__tmp99/loop ) );
    nor3_1 \cxe/Unr  ( .x(\cxe/nr ), .a(eop_ix), .b(nack_x), .c(sx) );
    nand3_1 \cxe/Und  ( .x(\cxe/nd ), .a(eop_ix), .b(nack_x), .c(sx) );
    oa21_1 \cxe/U1  ( .x(\cxe/n2 ), .a(\cxe/n2 ), .b(\cxe/nr ), .c(\cxe/nd )
         );
    inv_1 \cxe/U3  ( .x(eop_ox), .a(\cxe/n2 ) );
    ao31_1 \cx3/__tmp99/aoi  ( .x(\cx3/__tmp99/loop ), .a(d3_ix), .b(nack_x), 
        .c(sx), .d(d3_ox) );
    oa21_1 \cx3/__tmp99/outGate  ( .x(d3_ox), .a(d3_ix), .b(nack_x), .c(
        \cx3/__tmp99/loop ) );
    ao31_1 \cx2/__tmp99/aoi  ( .x(\cx2/__tmp99/loop ), .a(d2_ix), .b(nack_x), 
        .c(sx), .d(d2_ox) );
    oa21_1 \cx2/__tmp99/outGate  ( .x(d2_ox), .a(d2_ix), .b(nack_x), .c(
        \cx2/__tmp99/loop ) );
    ao31_1 \cx1/__tmp99/aoi  ( .x(\cx1/__tmp99/loop ), .a(d1_ix), .b(nack_x), 
        .c(sx), .d(d1_ox) );
    oa21_1 \cx1/__tmp99/outGate  ( .x(d1_ox), .a(d1_ix), .b(nack_x), .c(
        \cx1/__tmp99/loop ) );
    ao31_1 \cx0/__tmp99/aoi  ( .x(\cx0/__tmp99/loop ), .a(d0_ix), .b(nack_x), 
        .c(sx), .d(d0_ox) );
    oa21_1 \cx0/__tmp99/outGate  ( .x(d0_ox), .a(d0_ix), .b(nack_x), .c(
        \cx0/__tmp99/loop ) );
    nand2_1 \mtx/mg2  ( .x(\mtx/gr2 ), .a(mry), .b(\mtx/gr1 ) );
    nand2_1 \mtx/U1  ( .x(\mtx/gr1 ), .a(mrx), .b(\mtx/gr2 ) );
    nor3_1 \mtx/U2  ( .x(gy), .a(\mtx/gr2 ), .b(\mtx/gr2 ), .c(\mtx/gr2 ) );
    nor3_1 \mtx/U3  ( .x(gx), .a(\mtx/gr1 ), .b(\mtx/gr1 ), .c(\mtx/gr1 ) );
    nor2_1 \sry/i1  ( .x(\sry/qz ), .a(req_y), .b(mry) );
    nor2_1 \srx/i1  ( .x(\srx/qz ), .a(req_x), .b(mrx) );
    latn_1 \sl_sy/lph3  ( .q(sy), .d(\sl_sy/l1_q ), .g(phi3) );
    latn_1 \sl_sy/lph2  ( .q(\scan[1] ), .d(\sl_sy/l1_q ), .g(phi2) );
    mux2_1 \sl_sy/mxl/mux  ( .x(\sl_sy/mxl/muxout ), .d0(sy_pl), .sl(test_se), 
        .d1(\scan[0] ) );
    latn_1 \sl_sy/mxl/lph1  ( .q(\sl_sy/l1_q ), .d(\sl_sy/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_sx/lph3  ( .q(sx), .d(\sl_sx/l1_q ), .g(phi3) );
    latn_1 \sl_sx/lph2  ( .q(\scan[0] ), .d(\sl_sx/l1_q ), .g(phi2) );
    mux2_1 \sl_sx/mxl/mux  ( .x(\sl_sx/mxl/muxout ), .d0(sx_pl), .sl(test_se), 
        .d1(test_si) );
    latn_1 \sl_sx/mxl/lph1  ( .q(\sl_sx/l1_q ), .d(\sl_sx/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAcky/lph3  ( .q(acky_l), .d(\slAcky/l1_q ), .g(phi3) );
    latn_1 \slAcky/lph2  ( .q(test_so), .d(\slAcky/l1_q ), .g(phi2) );
    mux2_1 \slAcky/mxl/mux  ( .x(\slAcky/mxl/muxout ), .d0(ack_oxy), .sl(
        test_se), .d1(\scan[2] ) );
    latn_1 \slAcky/mxl/lph1  ( .q(\slAcky/l1_q ), .d(\slAcky/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAckx/lph3  ( .q(ackx_l), .d(\slAckx/l1_q ), .g(phi3) );
    latn_1 \slAckx/lph2  ( .q(\scan[2] ), .d(\slAckx/l1_q ), .g(phi2) );
    mux2_1 \slAckx/mxl/mux  ( .x(\slAckx/mxl/muxout ), .d0(ack_oxy), .sl(
        test_se), .d1(\scan[1] ) );
    latn_1 \slAckx/mxl/lph1  ( .q(\slAckx/l1_q ), .d(\slAckx/mxl/muxout ), .g(
        phi1) );
    nor3_1 U1 ( .x(mrx), .a(eop_ox), .b(rst), .c(\srx/qz ) );
    nor3_1 U2 ( .x(mry), .a(eop_oy), .b(rst), .c(\sry/qz ) );
endmodule


module chain_arbiter12 ( eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, ack_ix, eop_iy, 
    d0_iy, d1_iy, d2_iy, d3_iy, ack_iy, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, 
    eop_oy, d0_oy, d1_oy, d2_oy, d3_oy, ack_oxy, rst, test_si, test_se, 
    test_so, phi1, phi2, phi3 );
input  eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, eop_iy, d0_iy, d1_iy, d2_iy, d3_iy, 
    ack_oxy, rst, test_si, test_se, phi1, phi2, phi3;
output ack_ix, ack_iy, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, eop_oy, d0_oy, 
    d1_oy, d2_oy, d3_oy, test_so;
    wire \scan[1] , \scan[2] , ackx_l, nack_x, sx, acky_l, nack_y, sy, mrx, 
        req_x, mry, req_y, gx, gy, \scan[0] , sx_pl, sy_pl, n1x, n2x, n1y, n2y, 
        n5x, n6x, n5y, n6y, \cye/nr , \cye/nd , \cye/n2 , \cy3/__tmp99/loop , 
        \cy2/__tmp99/loop , \cy1/__tmp99/loop , \cy0/__tmp99/loop , \cxe/nr , 
        \cxe/nd , \cxe/n2 , \cx3/__tmp99/loop , \cx2/__tmp99/loop , 
        \cx1/__tmp99/loop , \cx0/__tmp99/loop , \mtx/gr2 , \mtx/gr1 , \sry/qz , 
        \srx/qz , \sl_sy/l1_q , \sl_sy/mxl/muxout , \sl_sx/l1_q , 
        \sl_sx/mxl/muxout , \slAcky/l1_q , \slAcky/mxl/muxout , \slAckx/l1_q , 
        \slAckx/mxl/muxout ;
    nor2_2 U12 ( .x(nack_x), .a(ackx_l), .b(rst) );
    nand2_1 U4 ( .x(ack_ix), .a(n1x), .b(n2x) );
    nor3_1 U17 ( .x(n1x), .a(d2_ox), .b(d3_ox), .c(d1_ox) );
    nor2_1 U18 ( .x(n2x), .a(eop_ox), .b(d0_ox) );
    nor2_2 U11 ( .x(nack_y), .a(acky_l), .b(rst) );
    nand2_1 U3 ( .x(ack_iy), .a(n1y), .b(n2y) );
    nor3_1 U16 ( .x(n1y), .a(d2_oy), .b(d3_oy), .c(d1_oy) );
    nor2_1 U19 ( .x(n2y), .a(eop_oy), .b(d0_oy) );
    nand2_1 U15 ( .x(req_x), .a(n5x), .b(n6x) );
    nor3_1 U10 ( .x(n5x), .a(d2_ix), .b(d3_ix), .c(d1_ix) );
    nor2_1 U13 ( .x(n6x), .a(eop_ix), .b(d0_ix) );
    nand2_1 U14 ( .x(req_y), .a(n5y), .b(n6y) );
    nor3_1 U9 ( .x(n5y), .a(d2_iy), .b(d3_iy), .c(d1_iy) );
    nor2_1 U20 ( .x(n6y), .a(eop_iy), .b(d0_iy) );
    nor2i_1 U6 ( .x(sx_pl), .a(gx), .b(eop_oy) );
    nor2i_1 U5 ( .x(sy_pl), .a(gy), .b(eop_ox) );
    nor3_1 \cye/Unr  ( .x(\cye/nr ), .a(eop_iy), .b(nack_y), .c(sy) );
    nand3_1 \cye/Und  ( .x(\cye/nd ), .a(eop_iy), .b(nack_y), .c(sy) );
    oa21_1 \cye/U1  ( .x(\cye/n2 ), .a(\cye/n2 ), .b(\cye/nr ), .c(\cye/nd )
         );
    inv_1 \cye/U3  ( .x(eop_oy), .a(\cye/n2 ) );
    ao31_1 \cy3/__tmp99/aoi  ( .x(\cy3/__tmp99/loop ), .a(d3_iy), .b(nack_y), 
        .c(sy), .d(d3_oy) );
    oa21_1 \cy3/__tmp99/outGate  ( .x(d3_oy), .a(d3_iy), .b(nack_y), .c(
        \cy3/__tmp99/loop ) );
    ao31_1 \cy2/__tmp99/aoi  ( .x(\cy2/__tmp99/loop ), .a(d2_iy), .b(nack_y), 
        .c(sy), .d(d2_oy) );
    oa21_1 \cy2/__tmp99/outGate  ( .x(d2_oy), .a(d2_iy), .b(nack_y), .c(
        \cy2/__tmp99/loop ) );
    ao31_1 \cy1/__tmp99/aoi  ( .x(\cy1/__tmp99/loop ), .a(d1_iy), .b(nack_y), 
        .c(sy), .d(d1_oy) );
    oa21_1 \cy1/__tmp99/outGate  ( .x(d1_oy), .a(d1_iy), .b(nack_y), .c(
        \cy1/__tmp99/loop ) );
    ao31_1 \cy0/__tmp99/aoi  ( .x(\cy0/__tmp99/loop ), .a(d0_iy), .b(nack_y), 
        .c(sy), .d(d0_oy) );
    oa21_1 \cy0/__tmp99/outGate  ( .x(d0_oy), .a(d0_iy), .b(nack_y), .c(
        \cy0/__tmp99/loop ) );
    nor3_1 \cxe/Unr  ( .x(\cxe/nr ), .a(eop_ix), .b(nack_x), .c(sx) );
    nand3_1 \cxe/Und  ( .x(\cxe/nd ), .a(eop_ix), .b(nack_x), .c(sx) );
    oa21_1 \cxe/U1  ( .x(\cxe/n2 ), .a(\cxe/n2 ), .b(\cxe/nr ), .c(\cxe/nd )
         );
    inv_1 \cxe/U3  ( .x(eop_ox), .a(\cxe/n2 ) );
    ao31_1 \cx3/__tmp99/aoi  ( .x(\cx3/__tmp99/loop ), .a(d3_ix), .b(nack_x), 
        .c(sx), .d(d3_ox) );
    oa21_1 \cx3/__tmp99/outGate  ( .x(d3_ox), .a(d3_ix), .b(nack_x), .c(
        \cx3/__tmp99/loop ) );
    ao31_1 \cx2/__tmp99/aoi  ( .x(\cx2/__tmp99/loop ), .a(d2_ix), .b(nack_x), 
        .c(sx), .d(d2_ox) );
    oa21_1 \cx2/__tmp99/outGate  ( .x(d2_ox), .a(d2_ix), .b(nack_x), .c(
        \cx2/__tmp99/loop ) );
    ao31_1 \cx1/__tmp99/aoi  ( .x(\cx1/__tmp99/loop ), .a(d1_ix), .b(nack_x), 
        .c(sx), .d(d1_ox) );
    oa21_1 \cx1/__tmp99/outGate  ( .x(d1_ox), .a(d1_ix), .b(nack_x), .c(
        \cx1/__tmp99/loop ) );
    ao31_1 \cx0/__tmp99/aoi  ( .x(\cx0/__tmp99/loop ), .a(d0_ix), .b(nack_x), 
        .c(sx), .d(d0_ox) );
    oa21_1 \cx0/__tmp99/outGate  ( .x(d0_ox), .a(d0_ix), .b(nack_x), .c(
        \cx0/__tmp99/loop ) );
    nand2_1 \mtx/mg2  ( .x(\mtx/gr2 ), .a(mry), .b(\mtx/gr1 ) );
    nand2_1 \mtx/U1  ( .x(\mtx/gr1 ), .a(mrx), .b(\mtx/gr2 ) );
    nor3_1 \mtx/U2  ( .x(gy), .a(\mtx/gr2 ), .b(\mtx/gr2 ), .c(\mtx/gr2 ) );
    nor3_1 \mtx/U3  ( .x(gx), .a(\mtx/gr1 ), .b(\mtx/gr1 ), .c(\mtx/gr1 ) );
    nor2_1 \sry/i1  ( .x(\sry/qz ), .a(req_y), .b(mry) );
    nor2_1 \srx/i1  ( .x(\srx/qz ), .a(req_x), .b(mrx) );
    latn_1 \sl_sy/lph3  ( .q(sy), .d(\sl_sy/l1_q ), .g(phi3) );
    latn_1 \sl_sy/lph2  ( .q(\scan[1] ), .d(\sl_sy/l1_q ), .g(phi2) );
    mux2_1 \sl_sy/mxl/mux  ( .x(\sl_sy/mxl/muxout ), .d0(sy_pl), .sl(test_se), 
        .d1(\scan[0] ) );
    latn_1 \sl_sy/mxl/lph1  ( .q(\sl_sy/l1_q ), .d(\sl_sy/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_sx/lph3  ( .q(sx), .d(\sl_sx/l1_q ), .g(phi3) );
    latn_1 \sl_sx/lph2  ( .q(\scan[0] ), .d(\sl_sx/l1_q ), .g(phi2) );
    mux2_1 \sl_sx/mxl/mux  ( .x(\sl_sx/mxl/muxout ), .d0(sx_pl), .sl(test_se), 
        .d1(test_si) );
    latn_1 \sl_sx/mxl/lph1  ( .q(\sl_sx/l1_q ), .d(\sl_sx/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAcky/lph3  ( .q(acky_l), .d(\slAcky/l1_q ), .g(phi3) );
    latn_1 \slAcky/lph2  ( .q(test_so), .d(\slAcky/l1_q ), .g(phi2) );
    mux2_1 \slAcky/mxl/mux  ( .x(\slAcky/mxl/muxout ), .d0(ack_oxy), .sl(
        test_se), .d1(\scan[2] ) );
    latn_1 \slAcky/mxl/lph1  ( .q(\slAcky/l1_q ), .d(\slAcky/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAckx/lph3  ( .q(ackx_l), .d(\slAckx/l1_q ), .g(phi3) );
    latn_1 \slAckx/lph2  ( .q(\scan[2] ), .d(\slAckx/l1_q ), .g(phi2) );
    mux2_1 \slAckx/mxl/mux  ( .x(\slAckx/mxl/muxout ), .d0(ack_oxy), .sl(
        test_se), .d1(\scan[1] ) );
    latn_1 \slAckx/mxl/lph1  ( .q(\slAckx/l1_q ), .d(\slAckx/mxl/muxout ), .g(
        phi1) );
    nor3_1 U1 ( .x(mry), .a(eop_oy), .b(rst), .c(\sry/qz ) );
    nor3_1 U2 ( .x(mrx), .a(eop_ox), .b(rst), .c(\srx/qz ) );
endmodule


module chain_mux10 ( eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, ack_ixy, eop_iy, 
    d0_iy, d1_iy, d2_iy, d3_iy, eop_o, d0_o, d1_o, d2_o, d3_o, ack_o, rst, 
    test_si, test_se, test_so, phi1, phi2, phi3 );
input  eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, eop_iy, d0_iy, d1_iy, d2_iy, d3_iy, 
    ack_o, rst, test_si, test_se, phi1, phi2, phi3;
output ack_ixy, eop_o, d0_o, d1_o, d2_o, d3_o, test_so;
    wire ack_l, d0_i, ack, d1_i, d2_i, d3_i, eop_i, n1, n2, \ce/ob , \c3/ob , 
        \c2/ob , \c1/ob , \c0/ob , \slAck/l1_q , \slAck/mxl/muxout ;
    nor2_1 U2 ( .x(d3_i), .a(d3_iy), .b(d3_ix) );
    nor2_1 U3 ( .x(d2_i), .a(d2_iy), .b(d2_ix) );
    nor2_1 U4 ( .x(d1_i), .a(d1_iy), .b(d1_ix) );
    nor2_1 U5 ( .x(d0_i), .a(d0_iy), .b(d0_ix) );
    nor2_1 U6 ( .x(eop_i), .a(eop_iy), .b(eop_ix) );
    nand2_1 U1 ( .x(ack_ixy), .a(n1), .b(n2) );
    nor3_1 U9 ( .x(n1), .a(d2_o), .b(d3_o), .c(d1_o) );
    nor2_1 U8 ( .x(n2), .a(eop_o), .b(d0_o) );
    inv_1 \ce/Ui  ( .x(\ce/ob ), .a(eop_o) );
    aoi222_1 \ce/__tmp99/U1  ( .x(eop_o), .a(eop_i), .b(ack), .c(eop_i), .d(
        \ce/ob ), .e(ack), .f(\ce/ob ) );
    inv_1 \c3/Ui  ( .x(\c3/ob ), .a(d3_o) );
    aoi222_1 \c3/__tmp99/U1  ( .x(d3_o), .a(d3_i), .b(ack), .c(d3_i), .d(
        \c3/ob ), .e(ack), .f(\c3/ob ) );
    inv_1 \c2/Ui  ( .x(\c2/ob ), .a(d2_o) );
    aoi222_1 \c2/__tmp99/U1  ( .x(d2_o), .a(d2_i), .b(ack), .c(d2_i), .d(
        \c2/ob ), .e(ack), .f(\c2/ob ) );
    inv_1 \c1/Ui  ( .x(\c1/ob ), .a(d1_o) );
    aoi222_1 \c1/__tmp99/U1  ( .x(d1_o), .a(d1_i), .b(ack), .c(d1_i), .d(
        \c1/ob ), .e(ack), .f(\c1/ob ) );
    inv_1 \c0/Ui  ( .x(\c0/ob ), .a(d0_o) );
    aoi222_1 \c0/__tmp99/U1  ( .x(d0_o), .a(d0_i), .b(ack), .c(d0_i), .d(
        \c0/ob ), .e(ack), .f(\c0/ob ) );
    latn_1 \slAck/lph3  ( .q(ack_l), .d(\slAck/l1_q ), .g(phi3) );
    latn_1 \slAck/lph2  ( .q(test_so), .d(\slAck/l1_q ), .g(phi2) );
    mux2_1 \slAck/mxl/mux  ( .x(\slAck/mxl/muxout ), .d0(ack_o), .sl(test_se), 
        .d1(test_si) );
    latn_1 \slAck/mxl/lph1  ( .q(\slAck/l1_q ), .d(\slAck/mxl/muxout ), .g(
        phi1) );
    or2_4 U7 ( .x(ack), .a(ack_l), .b(rst) );
endmodule


module chain_mux11 ( eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, ack_ixy, eop_iy, 
    d0_iy, d1_iy, d2_iy, d3_iy, eop_o, d0_o, d1_o, d2_o, d3_o, ack_o, rst, 
    test_si, test_se, test_so, phi1, phi2, phi3 );
input  eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, eop_iy, d0_iy, d1_iy, d2_iy, d3_iy, 
    ack_o, rst, test_si, test_se, phi1, phi2, phi3;
output ack_ixy, eop_o, d0_o, d1_o, d2_o, d3_o, test_so;
    wire ack_l, d0_i, ack, d1_i, d2_i, d3_i, eop_i, n1, n2, \ce/ob , \c3/ob , 
        \c2/ob , \c1/ob , \c0/ob , \slAck/l1_q , \slAck/mxl/muxout ;
    nor2_1 U2 ( .x(d3_i), .a(d3_iy), .b(d3_ix) );
    nor2_1 U3 ( .x(d2_i), .a(d2_iy), .b(d2_ix) );
    nor2_1 U4 ( .x(d1_i), .a(d1_iy), .b(d1_ix) );
    nor2_1 U5 ( .x(d0_i), .a(d0_iy), .b(d0_ix) );
    nor2_1 U6 ( .x(eop_i), .a(eop_iy), .b(eop_ix) );
    nand2_1 U1 ( .x(ack_ixy), .a(n1), .b(n2) );
    nor3_1 U9 ( .x(n1), .a(d2_o), .b(d3_o), .c(d1_o) );
    nor2_1 U8 ( .x(n2), .a(eop_o), .b(d0_o) );
    inv_1 \ce/Ui  ( .x(\ce/ob ), .a(eop_o) );
    aoi222_1 \ce/__tmp99/U1  ( .x(eop_o), .a(eop_i), .b(ack), .c(eop_i), .d(
        \ce/ob ), .e(ack), .f(\ce/ob ) );
    inv_1 \c3/Ui  ( .x(\c3/ob ), .a(d3_o) );
    aoi222_1 \c3/__tmp99/U1  ( .x(d3_o), .a(d3_i), .b(ack), .c(d3_i), .d(
        \c3/ob ), .e(ack), .f(\c3/ob ) );
    inv_1 \c2/Ui  ( .x(\c2/ob ), .a(d2_o) );
    aoi222_1 \c2/__tmp99/U1  ( .x(d2_o), .a(d2_i), .b(ack), .c(d2_i), .d(
        \c2/ob ), .e(ack), .f(\c2/ob ) );
    inv_1 \c1/Ui  ( .x(\c1/ob ), .a(d1_o) );
    aoi222_1 \c1/__tmp99/U1  ( .x(d1_o), .a(d1_i), .b(ack), .c(d1_i), .d(
        \c1/ob ), .e(ack), .f(\c1/ob ) );
    inv_1 \c0/Ui  ( .x(\c0/ob ), .a(d0_o) );
    aoi222_1 \c0/__tmp99/U1  ( .x(d0_o), .a(d0_i), .b(ack), .c(d0_i), .d(
        \c0/ob ), .e(ack), .f(\c0/ob ) );
    latn_1 \slAck/lph3  ( .q(ack_l), .d(\slAck/l1_q ), .g(phi3) );
    latn_1 \slAck/lph2  ( .q(test_so), .d(\slAck/l1_q ), .g(phi2) );
    mux2_1 \slAck/mxl/mux  ( .x(\slAck/mxl/muxout ), .d0(ack_o), .sl(test_se), 
        .d1(test_si) );
    latn_1 \slAck/mxl/lph1  ( .q(\slAck/l1_q ), .d(\slAck/mxl/muxout ), .g(
        phi1) );
    or2_4 U7 ( .x(ack), .a(ack_l), .b(rst) );
endmodule


module chain_mux12 ( eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, ack_ixy, eop_iy, 
    d0_iy, d1_iy, d2_iy, d3_iy, eop_o, d0_o, d1_o, d2_o, d3_o, ack_o, rst, 
    test_si, test_se, test_so, phi1, phi2, phi3 );
input  eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, eop_iy, d0_iy, d1_iy, d2_iy, d3_iy, 
    ack_o, rst, test_si, test_se, phi1, phi2, phi3;
output ack_ixy, eop_o, d0_o, d1_o, d2_o, d3_o, test_so;
    wire ack_l, d0_i, ack, d1_i, d2_i, d3_i, eop_i, n1, n2, \ce/ob , \c3/ob , 
        \c2/ob , \c1/ob , \c0/ob , \slAck/l1_q , \slAck/mxl/muxout ;
    nor2_1 U2 ( .x(d3_i), .a(d3_iy), .b(d3_ix) );
    nor2_1 U3 ( .x(d2_i), .a(d2_iy), .b(d2_ix) );
    nor2_1 U4 ( .x(d1_i), .a(d1_iy), .b(d1_ix) );
    nor2_1 U5 ( .x(d0_i), .a(d0_iy), .b(d0_ix) );
    nor2_1 U6 ( .x(eop_i), .a(eop_iy), .b(eop_ix) );
    nand2_1 U1 ( .x(ack_ixy), .a(n1), .b(n2) );
    nor3_1 U9 ( .x(n1), .a(d2_o), .b(d3_o), .c(d1_o) );
    nor2_1 U8 ( .x(n2), .a(eop_o), .b(d0_o) );
    inv_1 \ce/Ui  ( .x(\ce/ob ), .a(eop_o) );
    aoi222_1 \ce/__tmp99/U1  ( .x(eop_o), .a(eop_i), .b(ack), .c(eop_i), .d(
        \ce/ob ), .e(ack), .f(\ce/ob ) );
    inv_1 \c3/Ui  ( .x(\c3/ob ), .a(d3_o) );
    aoi222_1 \c3/__tmp99/U1  ( .x(d3_o), .a(d3_i), .b(ack), .c(d3_i), .d(
        \c3/ob ), .e(ack), .f(\c3/ob ) );
    inv_1 \c2/Ui  ( .x(\c2/ob ), .a(d2_o) );
    aoi222_1 \c2/__tmp99/U1  ( .x(d2_o), .a(d2_i), .b(ack), .c(d2_i), .d(
        \c2/ob ), .e(ack), .f(\c2/ob ) );
    inv_1 \c1/Ui  ( .x(\c1/ob ), .a(d1_o) );
    aoi222_1 \c1/__tmp99/U1  ( .x(d1_o), .a(d1_i), .b(ack), .c(d1_i), .d(
        \c1/ob ), .e(ack), .f(\c1/ob ) );
    inv_1 \c0/Ui  ( .x(\c0/ob ), .a(d0_o) );
    aoi222_1 \c0/__tmp99/U1  ( .x(d0_o), .a(d0_i), .b(ack), .c(d0_i), .d(
        \c0/ob ), .e(ack), .f(\c0/ob ) );
    latn_1 \slAck/lph3  ( .q(ack_l), .d(\slAck/l1_q ), .g(phi3) );
    latn_1 \slAck/lph2  ( .q(test_so), .d(\slAck/l1_q ), .g(phi2) );
    mux2_1 \slAck/mxl/mux  ( .x(\slAck/mxl/muxout ), .d0(ack_o), .sl(test_se), 
        .d1(test_si) );
    latn_1 \slAck/mxl/lph1  ( .q(\slAck/l1_q ), .d(\slAck/mxl/muxout ), .g(
        phi1) );
    or2_4 U7 ( .x(ack), .a(ack_l), .b(rst) );
endmodule


module resp_fab ( nrst, IMEM_eop_i, IMEM_d0_i, IMEM_d1_i, IMEM_d2_i, IMEM_d3_i, 
    IMEM_ack, DMEM_eop_i, DMEM_d0_i, DMEM_d1_i, DMEM_d2_i, DMEM_d3_i, DMEM_ack, 
    WB_eop_i, WB_d0_i, WB_d1_i, WB_d2_i, WB_d3_i, WB_ack, BC_eop_i, BC_d0_i, 
    BC_d1_i, BC_d2_i, BC_d3_i, BC_ack, I_port_eop_i, I_port_d0_i, I_port_d1_i, 
    I_port_d2_i, I_port_d3_i, I_port_ack, TIC_eop_i, TIC_d0_i, TIC_d1_i, 
    TIC_d2_i, TIC_d3_i, TIC_ack, D_port_eop_i, D_port_d0_i, D_port_d1_i, 
    D_port_d2_i, D_port_d3_i, D_port_ack, test_si, test_so, test_se, phi1, 
    phi2, phi3 );
input  nrst, IMEM_eop_i, IMEM_d0_i, IMEM_d1_i, IMEM_d2_i, IMEM_d3_i, 
    DMEM_eop_i, DMEM_d0_i, DMEM_d1_i, DMEM_d2_i, DMEM_d3_i, WB_eop_i, WB_d0_i, 
    WB_d1_i, WB_d2_i, WB_d3_i, BC_eop_i, BC_d0_i, BC_d1_i, BC_d2_i, BC_d3_i, 
    I_port_ack, TIC_ack, D_port_ack, test_si, test_se, phi1, phi2, phi3;
output IMEM_ack, DMEM_ack, WB_ack, BC_ack, I_port_eop_i, I_port_d0_i, 
    I_port_d1_i, I_port_d2_i, I_port_d3_i, TIC_eop_i, TIC_d0_i, TIC_d1_i, 
    TIC_d2_i, TIC_d3_i, D_port_eop_i, D_port_d0_i, D_port_d1_i, D_port_d2_i, 
    D_port_d3_i, test_so;
    wire A10_eop_o0, A10_d0_o0, A10_d1_o0, A10_d2_o0, A10_d3_o0, A10_eop_o1, 
        A10_d0_o1, A10_d1_o1, A10_d2_o1, A10_d3_o1, A10_ack, rst, \scan[7] , 
        \scan[6] , \scan[5] , \scan[4] , \scan[3] , \scan[2] , \scan[1] , 
        M10_eop, M10_d0, M10_d1, M10_d2, M10_d3, M10_ack, A11_eop_o0, 
        A11_d0_o0, A11_d1_o0, A11_d2_o0, A11_d3_o0, A11_eop_o1, A11_d0_o1, 
        A11_d1_o1, A11_d2_o1, A11_d3_o1, A11_ack, M11_eop, M11_d0, M11_d1, 
        M11_d2, M11_d3, M11_ack, A12_eop_o0, A12_d0_o0, A12_d1_o0, A12_d2_o0, 
        A12_d3_o0, A12_eop_o1, A12_d0_o1, A12_d1_o1, A12_d2_o1, A12_d3_o1, 
        A12_ack, M12_eop, M12_d0, M12_d1, M12_d2, M12_d3, M12_ack, R10_odd_eop, 
        R10_odd_d0, R10_odd_d1, R10_odd_d2, R10_odd_d3, R10_odd_ack, n1, n2, 
        n3, n4;
    chain_arbiter10 arb10 ( .eop_ix(IMEM_eop_i), .d0_ix(IMEM_d0_i), .d1_ix(
        IMEM_d1_i), .d2_ix(IMEM_d2_i), .d3_ix(IMEM_d3_i), .ack_ix(IMEM_ack), 
        .eop_iy(DMEM_eop_i), .d0_iy(DMEM_d0_i), .d1_iy(DMEM_d1_i), .d2_iy(
        DMEM_d2_i), .d3_iy(DMEM_d3_i), .ack_iy(DMEM_ack), .eop_ox(A10_eop_o0), 
        .d0_ox(A10_d0_o0), .d1_ox(A10_d1_o0), .d2_ox(A10_d2_o0), .d3_ox(
        A10_d3_o0), .eop_oy(A10_eop_o1), .d0_oy(A10_d0_o1), .d1_oy(A10_d1_o1), 
        .d2_oy(A10_d2_o1), .d3_oy(A10_d3_o1), .ack_oxy(A10_ack), .rst(rst), 
        .test_si(test_si), .test_se(test_se), .test_so(\scan[1] ), .phi1(phi1), 
        .phi2(phi2), .phi3(phi3) );
    chain_mux10 mux10 ( .eop_ix(A10_eop_o0), .d0_ix(A10_d0_o0), .d1_ix(
        A10_d1_o0), .d2_ix(A10_d2_o0), .d3_ix(A10_d3_o0), .ack_ixy(A10_ack), 
        .eop_iy(A10_eop_o1), .d0_iy(A10_d0_o1), .d1_iy(A10_d1_o1), .d2_iy(
        A10_d2_o1), .d3_iy(A10_d3_o1), .eop_o(M10_eop), .d0_o(M10_d0), .d1_o(
        M10_d1), .d2_o(M10_d2), .d3_o(M10_d3), .ack_o(M10_ack), .rst(rst), 
        .test_si(\scan[1] ), .test_se(n4), .test_so(\scan[2] ), .phi1(n2), 
        .phi2(n1), .phi3(n3) );
    chain_arbiter11 arb11 ( .eop_ix(M10_eop), .d0_ix(M10_d0), .d1_ix(M10_d1), 
        .d2_ix(M10_d2), .d3_ix(M10_d3), .ack_ix(M10_ack), .eop_iy(BC_eop_i), 
        .d0_iy(BC_d0_i), .d1_iy(BC_d1_i), .d2_iy(BC_d2_i), .d3_iy(BC_d3_i), 
        .ack_iy(BC_ack), .eop_ox(A11_eop_o0), .d0_ox(A11_d0_o0), .d1_ox(
        A11_d1_o0), .d2_ox(A11_d2_o0), .d3_ox(A11_d3_o0), .eop_oy(A11_eop_o1), 
        .d0_oy(A11_d0_o1), .d1_oy(A11_d1_o1), .d2_oy(A11_d2_o1), .d3_oy(
        A11_d3_o1), .ack_oxy(A11_ack), .rst(rst), .test_si(\scan[2] ), 
        .test_se(n4), .test_so(\scan[3] ), .phi1(n2), .phi2(n1), .phi3(n3) );
    chain_mux11 mux11 ( .eop_ix(A11_eop_o0), .d0_ix(A11_d0_o0), .d1_ix(
        A11_d1_o0), .d2_ix(A11_d2_o0), .d3_ix(A11_d3_o0), .ack_ixy(A11_ack), 
        .eop_iy(A11_eop_o1), .d0_iy(A11_d0_o1), .d1_iy(A11_d1_o1), .d2_iy(
        A11_d2_o1), .d3_iy(A11_d3_o1), .eop_o(M11_eop), .d0_o(M11_d0), .d1_o(
        M11_d1), .d2_o(M11_d2), .d3_o(M11_d3), .ack_o(M11_ack), .rst(rst), 
        .test_si(\scan[3] ), .test_se(test_se), .test_so(\scan[4] ), .phi1(
        phi1), .phi2(phi2), .phi3(phi3) );
    chain_arbiter12 arb12 ( .eop_ix(M11_eop), .d0_ix(M11_d0), .d1_ix(M11_d1), 
        .d2_ix(M11_d2), .d3_ix(M11_d3), .ack_ix(M11_ack), .eop_iy(WB_eop_i), 
        .d0_iy(WB_d0_i), .d1_iy(WB_d1_i), .d2_iy(WB_d2_i), .d3_iy(WB_d3_i), 
        .ack_iy(WB_ack), .eop_ox(A12_eop_o0), .d0_ox(A12_d0_o0), .d1_ox(
        A12_d1_o0), .d2_ox(A12_d2_o0), .d3_ox(A12_d3_o0), .eop_oy(A12_eop_o1), 
        .d0_oy(A12_d0_o1), .d1_oy(A12_d1_o1), .d2_oy(A12_d2_o1), .d3_oy(
        A12_d3_o1), .ack_oxy(A12_ack), .rst(rst), .test_si(\scan[4] ), 
        .test_se(n4), .test_so(\scan[5] ), .phi1(n2), .phi2(n1), .phi3(n3) );
    chain_mux12 mux12 ( .eop_ix(A12_eop_o0), .d0_ix(A12_d0_o0), .d1_ix(
        A12_d1_o0), .d2_ix(A12_d2_o0), .d3_ix(A12_d3_o0), .ack_ixy(A12_ack), 
        .eop_iy(A12_eop_o1), .d0_iy(A12_d0_o1), .d1_iy(A12_d1_o1), .d2_iy(
        A12_d2_o1), .d3_iy(A12_d3_o1), .eop_o(M12_eop), .d0_o(M12_d0), .d1_o(
        M12_d1), .d2_o(M12_d2), .d3_o(M12_d3), .ack_o(M12_ack), .rst(rst), 
        .test_si(\scan[5] ), .test_se(n4), .test_so(\scan[6] ), .phi1(n2), 
        .phi2(n1), .phi3(n3) );
    chain_router10 router10 ( .eop_i(M12_eop), .d0_i(M12_d0), .d1_i(M12_d1), 
        .d2_i(M12_d2), .d3_i(M12_d3), .ack_i(M12_ack), .eop_ox(R10_odd_eop), 
        .d0_ox(R10_odd_d0), .d1_ox(R10_odd_d1), .d2_ox(R10_odd_d2), .d3_ox(
        R10_odd_d3), .ack_ox(R10_odd_ack), .eop_oy(TIC_eop_i), .d0_oy(TIC_d0_i
        ), .d1_oy(TIC_d1_i), .d2_oy(TIC_d2_i), .d3_oy(TIC_d3_i), .ack_oy(
        TIC_ack), .nrst(nrst), .test_si(\scan[6] ), .test_se(n4), .test_so(
        \scan[7] ), .phi1(phi1), .phi2(phi2), .phi3(phi3) );
    chain_router11 router11 ( .eop_i(R10_odd_eop), .d0_i(R10_odd_d0), .d1_i(
        R10_odd_d1), .d2_i(R10_odd_d2), .d3_i(R10_odd_d3), .ack_i(R10_odd_ack), 
        .eop_ox(I_port_eop_i), .d0_ox(I_port_d0_i), .d1_ox(I_port_d1_i), 
        .d2_ox(I_port_d2_i), .d3_ox(I_port_d3_i), .ack_ox(I_port_ack), 
        .eop_oy(D_port_eop_i), .d0_oy(D_port_d0_i), .d1_oy(D_port_d1_i), 
        .d2_oy(D_port_d2_i), .d3_oy(D_port_d3_i), .ack_oy(D_port_ack), .nrst(
        nrst), .test_si(\scan[7] ), .test_se(test_se), .test_so(test_so), 
        .phi1(phi1), .phi2(phi2), .phi3(phi3) );
    buf_1 U1 ( .x(n1), .a(phi2) );
    buf_1 U2 ( .x(n2), .a(phi1) );
    buf_1 U3 ( .x(n3), .a(phi3) );
    buf_3 U4 ( .x(n4), .a(test_se) );
    inv_5 U5 ( .x(rst), .a(nrst) );
endmodule


module resp_fab_scan ( nrst, IMEM_eop_i, IMEM_d0_i, IMEM_d1_i, IMEM_d2_i, 
    IMEM_d3_i, IMEM_ack, DMEM_eop_i, DMEM_d0_i, DMEM_d1_i, DMEM_d2_i, 
    DMEM_d3_i, DMEM_ack, WB_eop_i, WB_d0_i, WB_d1_i, WB_d2_i, WB_d3_i, WB_ack, 
    BC_eop_i, BC_d0_i, BC_d1_i, BC_d2_i, BC_d3_i, BC_ack, I_port_eop_i, 
    I_port_d0_i, I_port_d1_i, I_port_d2_i, I_port_d3_i, I_port_ack, TIC_eop_i, 
    TIC_d0_i, TIC_d1_i, TIC_d2_i, TIC_d3_i, TIC_ack, D_port_eop_i, D_port_d0_i, 
    D_port_d1_i, D_port_d2_i, D_port_d3_i, D_port_ack, test_si, test_so, 
    test_se, phi1, phi2, phi3 );
input  nrst, IMEM_eop_i, IMEM_d0_i, IMEM_d1_i, IMEM_d2_i, IMEM_d3_i, 
    DMEM_eop_i, DMEM_d0_i, DMEM_d1_i, DMEM_d2_i, DMEM_d3_i, WB_eop_i, WB_d0_i, 
    WB_d1_i, WB_d2_i, WB_d3_i, BC_eop_i, BC_d0_i, BC_d1_i, BC_d2_i, BC_d3_i, 
    I_port_ack, TIC_ack, D_port_ack, test_si, test_se, phi1, phi2, phi3;
output IMEM_ack, DMEM_ack, WB_ack, BC_ack, I_port_eop_i, I_port_d0_i, 
    I_port_d1_i, I_port_d2_i, I_port_d3_i, TIC_eop_i, TIC_d0_i, TIC_d1_i, 
    TIC_d2_i, TIC_d3_i, D_port_eop_i, D_port_d0_i, D_port_d1_i, D_port_d2_i, 
    D_port_d3_i, test_so;
    wire \scan[12] , \scan[11] , \scan[10] , \scan[9] , \scan[8] , \scan[7] , 
        \scan[6] , \scan[5] , \scan[4] , \scan[3] , \scan[2] , \scan[1] , 
        IMEM_eop_i_sc, IMEM_d0_i_sc, IMEM_d1_i_sc, IMEM_d2_i_sc, IMEM_d3_i_sc, 
        DMEM_eop_i_sc, DMEM_d0_i_sc, DMEM_d1_i_sc, DMEM_d2_i_sc, DMEM_d3_i_sc, 
        WB_eop_i_sc, WB_d0_i_sc, WB_d1_i_sc, WB_d2_i_sc, WB_d3_i_sc, 
        I_port_ack_sc, TIC_ack_sc, D_port_ack_sc, scan_m10, scan_m11, scan_m12, 
        \sc12_m_wbAck/muxout , \sc11_m_dmAck/muxout , \sc10_m_imAck/muxout , 
        \sc6_dpAck/l1_q , \sc6_dpAck/mxl/muxout , \sc5_ticAck/l1_q , 
        \sc5_ticAck/mxl/muxout , \sc4_ipAck/l1_q , \sc4_ipAck/mxl/muxout , 
        \sc_dp/intI0 , \sc_dp/scn0 , \sc_dp/intI1 , \sc_dp/scn1 , 
        \sc_dp/intI2 , \sc_dp/scn2 , \sc_dp/intI3 , \sc_dp/scn3 , 
        \sc_dp/intI4 , \sc_dp/l4_m/muxout , \sc_dp/l3_m/muxout , 
        \sc_dp/l2_m/muxout , \sc_dp/l1_m/muxout , \sc_dp/l0_m/muxout , 
        \sc_tic/intI0 , \sc_tic/scn0 , \sc_tic/intI1 , \sc_tic/scn1 , 
        \sc_tic/intI2 , \sc_tic/scn2 , \sc_tic/intI3 , \sc_tic/scn3 , 
        \sc_tic/intI4 , \sc_tic/l4_m/muxout , \sc_tic/l3_m/muxout , 
        \sc_tic/l2_m/muxout , \sc_tic/l1_m/muxout , \sc_tic/l0_m/muxout , 
        \sc_ip/intI0 , \sc_ip/scn0 , \sc_ip/intI1 , \sc_ip/scn1 , 
        \sc_ip/intI2 , \sc_ip/scn2 , \sc_ip/intI3 , \sc_ip/scn3 , 
        \sc_ip/intI4 , \sc_ip/l4_m/muxout , \sc_ip/l3_m/muxout , 
        \sc_ip/l2_m/muxout , \sc_ip/l1_m/muxout , \sc_ip/l0_m/muxout , 
        \sc_wb/scn1 , \sc_wb/scn2 , \sc_wb/scn3 , \sc_wb/scn4 , 
        \sc_wb/sl4/l1_q , \sc_wb/sl4/mxl/muxout , \sc_wb/sl3/l1_q , 
        \sc_wb/sl3/mxl/muxout , \sc_wb/sl2/l1_q , \sc_wb/sl2/mxl/muxout , 
        \sc_wb/sl1/l1_q , \sc_wb/sl1/mxl/muxout , \sc_wb/sl0/l1_q , 
        \sc_wb/sl0/mxl/muxout , \sc_dm/scn1 , \sc_dm/scn2 , \sc_dm/scn3 , 
        \sc_dm/scn4 , \sc_dm/sl4/l1_q , \sc_dm/sl4/mxl/muxout , 
        \sc_dm/sl3/l1_q , \sc_dm/sl3/mxl/muxout , \sc_dm/sl2/l1_q , 
        \sc_dm/sl2/mxl/muxout , \sc_dm/sl1/l1_q , \sc_dm/sl1/mxl/muxout , 
        \sc_dm/sl0/l1_q , \sc_dm/sl0/mxl/muxout , \sc_im/scn1 , \sc_im/scn2 , 
        \sc_im/scn3 , \sc_im/scn4 , \sc_im/sl4/l1_q , \sc_im/sl4/mxl/muxout , 
        \sc_im/sl3/l1_q , \sc_im/sl3/mxl/muxout , \sc_im/sl2/l1_q , 
        \sc_im/sl2/mxl/muxout , \sc_im/sl1/l1_q , \sc_im/sl1/mxl/muxout , 
        \sc_im/sl0/l1_q , \sc_im/sl0/mxl/muxout , n1, n2, n3, n4, n5, n6, n7, 
        n8, n9, n10, n11, n12, n13, n14, n15;
    resp_fab fab2 ( .nrst(nrst), .IMEM_eop_i(IMEM_eop_i_sc), .IMEM_d0_i(
        IMEM_d0_i_sc), .IMEM_d1_i(IMEM_d1_i_sc), .IMEM_d2_i(IMEM_d2_i_sc), 
        .IMEM_d3_i(IMEM_d3_i_sc), .IMEM_ack(IMEM_ack), .DMEM_eop_i(
        DMEM_eop_i_sc), .DMEM_d0_i(DMEM_d0_i_sc), .DMEM_d1_i(DMEM_d1_i_sc), 
        .DMEM_d2_i(DMEM_d2_i_sc), .DMEM_d3_i(DMEM_d3_i_sc), .DMEM_ack(DMEM_ack
        ), .WB_eop_i(WB_eop_i_sc), .WB_d0_i(WB_d0_i_sc), .WB_d1_i(WB_d1_i_sc), 
        .WB_d2_i(WB_d2_i_sc), .WB_d3_i(WB_d3_i_sc), .WB_ack(WB_ack), 
        .BC_eop_i(BC_eop_i), .BC_d0_i(BC_d0_i), .BC_d1_i(BC_d1_i), .BC_d2_i(
        BC_d2_i), .BC_d3_i(BC_d3_i), .BC_ack(BC_ack), .I_port_eop_i(
        I_port_eop_i), .I_port_d0_i(I_port_d0_i), .I_port_d1_i(I_port_d1_i), 
        .I_port_d2_i(I_port_d2_i), .I_port_d3_i(I_port_d3_i), .I_port_ack(
        I_port_ack_sc), .TIC_eop_i(TIC_eop_i), .TIC_d0_i(TIC_d0_i), .TIC_d1_i(
        TIC_d1_i), .TIC_d2_i(TIC_d2_i), .TIC_d3_i(TIC_d3_i), .TIC_ack(
        TIC_ack_sc), .D_port_eop_i(D_port_eop_i), .D_port_d0_i(D_port_d0_i), 
        .D_port_d1_i(D_port_d1_i), .D_port_d2_i(D_port_d2_i), .D_port_d3_i(
        D_port_d3_i), .D_port_ack(D_port_ack_sc), .test_si(\scan[6] ), 
        .test_so(\scan[7] ), .test_se(n5), .phi1(n9), .phi2(n13), .phi3(n2) );
    latn_1 sc10_s_imAck ( .q(\scan[11] ), .d(scan_m10), .g(n15) );
    latn_1 sc11_s_dmAck ( .q(\scan[12] ), .d(scan_m11), .g(n12) );
    latn_1 sc12_s_wbAck ( .q(test_so), .d(scan_m12), .g(n14) );
    mux2_1 \sc12_m_wbAck/mux  ( .x(\sc12_m_wbAck/muxout ), .d0(WB_ack), .sl(n7
        ), .d1(\scan[12] ) );
    latn_1 \sc12_m_wbAck/lph1  ( .q(scan_m12), .d(\sc12_m_wbAck/muxout ), .g(
        n11) );
    mux2_1 \sc11_m_dmAck/mux  ( .x(\sc11_m_dmAck/muxout ), .d0(DMEM_ack), .sl(
        n6), .d1(\scan[11] ) );
    latn_1 \sc11_m_dmAck/lph1  ( .q(scan_m11), .d(\sc11_m_dmAck/muxout ), .g(
        n8) );
    mux2_1 \sc10_m_imAck/mux  ( .x(\sc10_m_imAck/muxout ), .d0(IMEM_ack), .sl(
        n6), .d1(\scan[10] ) );
    latn_1 \sc10_m_imAck/lph1  ( .q(scan_m10), .d(\sc10_m_imAck/muxout ), .g(
        n10) );
    latn_1 \sc6_dpAck/lph3  ( .q(D_port_ack_sc), .d(\sc6_dpAck/l1_q ), .g(n1)
         );
    latn_1 \sc6_dpAck/lph2  ( .q(\scan[6] ), .d(\sc6_dpAck/l1_q ), .g(n15) );
    mux2_1 \sc6_dpAck/mxl/mux  ( .x(\sc6_dpAck/mxl/muxout ), .d0(D_port_ack), 
        .sl(n7), .d1(\scan[5] ) );
    latn_1 \sc6_dpAck/mxl/lph1  ( .q(\sc6_dpAck/l1_q ), .d(
        \sc6_dpAck/mxl/muxout ), .g(n10) );
    latn_1 \sc5_ticAck/lph3  ( .q(TIC_ack_sc), .d(\sc5_ticAck/l1_q ), .g(n1)
         );
    latn_1 \sc5_ticAck/lph2  ( .q(\scan[5] ), .d(\sc5_ticAck/l1_q ), .g(n12)
         );
    mux2_1 \sc5_ticAck/mxl/mux  ( .x(\sc5_ticAck/mxl/muxout ), .d0(TIC_ack), 
        .sl(n4), .d1(\scan[4] ) );
    latn_1 \sc5_ticAck/mxl/lph1  ( .q(\sc5_ticAck/l1_q ), .d(
        \sc5_ticAck/mxl/muxout ), .g(n8) );
    latn_1 \sc4_ipAck/lph3  ( .q(I_port_ack_sc), .d(\sc4_ipAck/l1_q ), .g(n1)
         );
    latn_1 \sc4_ipAck/lph2  ( .q(\scan[4] ), .d(\sc4_ipAck/l1_q ), .g(n14) );
    mux2_1 \sc4_ipAck/mxl/mux  ( .x(\sc4_ipAck/mxl/muxout ), .d0(I_port_ack), 
        .sl(n4), .d1(\scan[3] ) );
    latn_1 \sc4_ipAck/mxl/lph1  ( .q(\sc4_ipAck/l1_q ), .d(
        \sc4_ipAck/mxl/muxout ), .g(n11) );
    latn_1 \sc_dp/l4_s  ( .q(\scan[10] ), .d(\sc_dp/intI4 ), .g(n15) );
    latn_1 \sc_dp/l3_s  ( .q(\sc_dp/scn3 ), .d(\sc_dp/intI3 ), .g(n12) );
    latn_1 \sc_dp/l2_s  ( .q(\sc_dp/scn2 ), .d(\sc_dp/intI2 ), .g(n14) );
    latn_1 \sc_dp/l1_s  ( .q(\sc_dp/scn1 ), .d(\sc_dp/intI1 ), .g(n15) );
    latn_1 \sc_dp/l0_s  ( .q(\sc_dp/scn0 ), .d(\sc_dp/intI0 ), .g(n12) );
    mux2_1 \sc_dp/l4_m/mux  ( .x(\sc_dp/l4_m/muxout ), .d0(D_port_d3_i), .sl(
        n4), .d1(\sc_dp/scn3 ) );
    latn_1 \sc_dp/l4_m/lph1  ( .q(\sc_dp/intI4 ), .d(\sc_dp/l4_m/muxout ), .g(
        n8) );
    mux2_1 \sc_dp/l3_m/mux  ( .x(\sc_dp/l3_m/muxout ), .d0(D_port_d2_i), .sl(
        n7), .d1(\sc_dp/scn2 ) );
    latn_1 \sc_dp/l3_m/lph1  ( .q(\sc_dp/intI3 ), .d(\sc_dp/l3_m/muxout ), .g(
        n11) );
    mux2_1 \sc_dp/l2_m/mux  ( .x(\sc_dp/l2_m/muxout ), .d0(D_port_d1_i), .sl(
        n6), .d1(\sc_dp/scn1 ) );
    latn_1 \sc_dp/l2_m/lph1  ( .q(\sc_dp/intI2 ), .d(\sc_dp/l2_m/muxout ), .g(
        n10) );
    mux2_1 \sc_dp/l1_m/mux  ( .x(\sc_dp/l1_m/muxout ), .d0(D_port_d0_i), .sl(
        n4), .d1(\sc_dp/scn0 ) );
    latn_1 \sc_dp/l1_m/lph1  ( .q(\sc_dp/intI1 ), .d(\sc_dp/l1_m/muxout ), .g(
        n8) );
    mux2_1 \sc_dp/l0_m/mux  ( .x(\sc_dp/l0_m/muxout ), .d0(D_port_eop_i), .sl(
        n7), .d1(\scan[9] ) );
    latn_1 \sc_dp/l0_m/lph1  ( .q(\sc_dp/intI0 ), .d(\sc_dp/l0_m/muxout ), .g(
        n11) );
    latn_1 \sc_tic/l4_s  ( .q(\scan[9] ), .d(\sc_tic/intI4 ), .g(n12) );
    latn_1 \sc_tic/l3_s  ( .q(\sc_tic/scn3 ), .d(\sc_tic/intI3 ), .g(n14) );
    latn_1 \sc_tic/l2_s  ( .q(\sc_tic/scn2 ), .d(\sc_tic/intI2 ), .g(n15) );
    latn_1 \sc_tic/l1_s  ( .q(\sc_tic/scn1 ), .d(\sc_tic/intI1 ), .g(n12) );
    latn_1 \sc_tic/l0_s  ( .q(\sc_tic/scn0 ), .d(\sc_tic/intI0 ), .g(n14) );
    mux2_1 \sc_tic/l4_m/mux  ( .x(\sc_tic/l4_m/muxout ), .d0(TIC_d3_i), .sl(n6
        ), .d1(\sc_tic/scn3 ) );
    latn_1 \sc_tic/l4_m/lph1  ( .q(\sc_tic/intI4 ), .d(\sc_tic/l4_m/muxout ), 
        .g(n10) );
    mux2_1 \sc_tic/l3_m/mux  ( .x(\sc_tic/l3_m/muxout ), .d0(TIC_d2_i), .sl(n4
        ), .d1(\sc_tic/scn2 ) );
    latn_1 \sc_tic/l3_m/lph1  ( .q(\sc_tic/intI3 ), .d(\sc_tic/l3_m/muxout ), 
        .g(n8) );
    mux2_1 \sc_tic/l2_m/mux  ( .x(\sc_tic/l2_m/muxout ), .d0(TIC_d1_i), .sl(n7
        ), .d1(\sc_tic/scn1 ) );
    latn_1 \sc_tic/l2_m/lph1  ( .q(\sc_tic/intI2 ), .d(\sc_tic/l2_m/muxout ), 
        .g(n11) );
    mux2_1 \sc_tic/l1_m/mux  ( .x(\sc_tic/l1_m/muxout ), .d0(TIC_d0_i), .sl(n6
        ), .d1(\sc_tic/scn0 ) );
    latn_1 \sc_tic/l1_m/lph1  ( .q(\sc_tic/intI1 ), .d(\sc_tic/l1_m/muxout ), 
        .g(n10) );
    mux2_1 \sc_tic/l0_m/mux  ( .x(\sc_tic/l0_m/muxout ), .d0(TIC_eop_i), .sl(
        n4), .d1(\scan[8] ) );
    latn_1 \sc_tic/l0_m/lph1  ( .q(\sc_tic/intI0 ), .d(\sc_tic/l0_m/muxout ), 
        .g(n8) );
    latn_1 \sc_ip/l4_s  ( .q(\scan[8] ), .d(\sc_ip/intI4 ), .g(n14) );
    latn_1 \sc_ip/l3_s  ( .q(\sc_ip/scn3 ), .d(\sc_ip/intI3 ), .g(n15) );
    latn_1 \sc_ip/l2_s  ( .q(\sc_ip/scn2 ), .d(\sc_ip/intI2 ), .g(n12) );
    latn_1 \sc_ip/l1_s  ( .q(\sc_ip/scn1 ), .d(\sc_ip/intI1 ), .g(n14) );
    latn_1 \sc_ip/l0_s  ( .q(\sc_ip/scn0 ), .d(\sc_ip/intI0 ), .g(n15) );
    mux2_1 \sc_ip/l4_m/mux  ( .x(\sc_ip/l4_m/muxout ), .d0(I_port_d3_i), .sl(
        n7), .d1(\sc_ip/scn3 ) );
    latn_1 \sc_ip/l4_m/lph1  ( .q(\sc_ip/intI4 ), .d(\sc_ip/l4_m/muxout ), .g(
        n11) );
    mux2_1 \sc_ip/l3_m/mux  ( .x(\sc_ip/l3_m/muxout ), .d0(I_port_d2_i), .sl(
        n7), .d1(\sc_ip/scn2 ) );
    latn_1 \sc_ip/l3_m/lph1  ( .q(\sc_ip/intI3 ), .d(\sc_ip/l3_m/muxout ), .g(
        n10) );
    mux2_1 \sc_ip/l2_m/mux  ( .x(\sc_ip/l2_m/muxout ), .d0(I_port_d1_i), .sl(
        n6), .d1(\sc_ip/scn1 ) );
    latn_1 \sc_ip/l2_m/lph1  ( .q(\sc_ip/intI2 ), .d(\sc_ip/l2_m/muxout ), .g(
        n8) );
    mux2_1 \sc_ip/l1_m/mux  ( .x(\sc_ip/l1_m/muxout ), .d0(I_port_d0_i), .sl(
        n4), .d1(\sc_ip/scn0 ) );
    latn_1 \sc_ip/l1_m/lph1  ( .q(\sc_ip/intI1 ), .d(\sc_ip/l1_m/muxout ), .g(
        n11) );
    mux2_1 \sc_ip/l0_m/mux  ( .x(\sc_ip/l0_m/muxout ), .d0(I_port_eop_i), .sl(
        n7), .d1(\scan[7] ) );
    latn_1 \sc_ip/l0_m/lph1  ( .q(\sc_ip/intI0 ), .d(\sc_ip/l0_m/muxout ), .g(
        n10) );
    latn_1 \sc_wb/sl4/lph3  ( .q(WB_d3_i_sc), .d(\sc_wb/sl4/l1_q ), .g(n3) );
    latn_1 \sc_wb/sl4/lph2  ( .q(\scan[3] ), .d(\sc_wb/sl4/l1_q ), .g(n12) );
    mux2_1 \sc_wb/sl4/mxl/mux  ( .x(\sc_wb/sl4/mxl/muxout ), .d0(WB_d3_i), 
        .sl(n6), .d1(\sc_wb/scn4 ) );
    latn_1 \sc_wb/sl4/mxl/lph1  ( .q(\sc_wb/sl4/l1_q ), .d(
        \sc_wb/sl4/mxl/muxout ), .g(n8) );
    latn_1 \sc_wb/sl3/lph3  ( .q(WB_d2_i_sc), .d(\sc_wb/sl3/l1_q ), .g(n3) );
    latn_1 \sc_wb/sl3/lph2  ( .q(\sc_wb/scn4 ), .d(\sc_wb/sl3/l1_q ), .g(n15)
         );
    mux2_1 \sc_wb/sl3/mxl/mux  ( .x(\sc_wb/sl3/mxl/muxout ), .d0(WB_d2_i), 
        .sl(n4), .d1(\sc_wb/scn3 ) );
    latn_1 \sc_wb/sl3/mxl/lph1  ( .q(\sc_wb/sl3/l1_q ), .d(
        \sc_wb/sl3/mxl/muxout ), .g(n11) );
    latn_1 \sc_wb/sl2/lph3  ( .q(WB_d1_i_sc), .d(\sc_wb/sl2/l1_q ), .g(n3) );
    latn_1 \sc_wb/sl2/lph2  ( .q(\sc_wb/scn3 ), .d(\sc_wb/sl2/l1_q ), .g(n14)
         );
    mux2_1 \sc_wb/sl2/mxl/mux  ( .x(\sc_wb/sl2/mxl/muxout ), .d0(WB_d1_i), 
        .sl(n7), .d1(\sc_wb/scn2 ) );
    latn_1 \sc_wb/sl2/mxl/lph1  ( .q(\sc_wb/sl2/l1_q ), .d(
        \sc_wb/sl2/mxl/muxout ), .g(n10) );
    latn_1 \sc_wb/sl1/lph3  ( .q(WB_d0_i_sc), .d(\sc_wb/sl1/l1_q ), .g(n3) );
    latn_1 \sc_wb/sl1/lph2  ( .q(\sc_wb/scn2 ), .d(\sc_wb/sl1/l1_q ), .g(n15)
         );
    mux2_1 \sc_wb/sl1/mxl/mux  ( .x(\sc_wb/sl1/mxl/muxout ), .d0(WB_d0_i), 
        .sl(n4), .d1(\sc_wb/scn1 ) );
    latn_1 \sc_wb/sl1/mxl/lph1  ( .q(\sc_wb/sl1/l1_q ), .d(
        \sc_wb/sl1/mxl/muxout ), .g(n11) );
    latn_1 \sc_wb/sl0/lph3  ( .q(WB_eop_i_sc), .d(\sc_wb/sl0/l1_q ), .g(n3) );
    latn_1 \sc_wb/sl0/lph2  ( .q(\sc_wb/scn1 ), .d(\sc_wb/sl0/l1_q ), .g(n12)
         );
    mux2_1 \sc_wb/sl0/mxl/mux  ( .x(\sc_wb/sl0/mxl/muxout ), .d0(WB_eop_i), 
        .sl(n4), .d1(\scan[2] ) );
    latn_1 \sc_wb/sl0/mxl/lph1  ( .q(\sc_wb/sl0/l1_q ), .d(
        \sc_wb/sl0/mxl/muxout ), .g(n8) );
    latn_1 \sc_dm/sl4/lph3  ( .q(DMEM_d3_i_sc), .d(\sc_dm/sl4/l1_q ), .g(n3)
         );
    latn_1 \sc_dm/sl4/lph2  ( .q(\scan[2] ), .d(\sc_dm/sl4/l1_q ), .g(n14) );
    mux2_1 \sc_dm/sl4/mxl/mux  ( .x(\sc_dm/sl4/mxl/muxout ), .d0(DMEM_d3_i), 
        .sl(n6), .d1(\sc_dm/scn4 ) );
    latn_1 \sc_dm/sl4/mxl/lph1  ( .q(\sc_dm/sl4/l1_q ), .d(
        \sc_dm/sl4/mxl/muxout ), .g(n10) );
    latn_1 \sc_dm/sl3/lph3  ( .q(DMEM_d2_i_sc), .d(\sc_dm/sl3/l1_q ), .g(n3)
         );
    latn_1 \sc_dm/sl3/lph2  ( .q(\sc_dm/scn4 ), .d(\sc_dm/sl3/l1_q ), .g(n15)
         );
    mux2_1 \sc_dm/sl3/mxl/mux  ( .x(\sc_dm/sl3/mxl/muxout ), .d0(DMEM_d2_i), 
        .sl(n7), .d1(\sc_dm/scn3 ) );
    latn_1 \sc_dm/sl3/mxl/lph1  ( .q(\sc_dm/sl3/l1_q ), .d(
        \sc_dm/sl3/mxl/muxout ), .g(n11) );
    latn_1 \sc_dm/sl2/lph3  ( .q(DMEM_d1_i_sc), .d(\sc_dm/sl2/l1_q ), .g(n3)
         );
    latn_1 \sc_dm/sl2/lph2  ( .q(\sc_dm/scn3 ), .d(\sc_dm/sl2/l1_q ), .g(n12)
         );
    mux2_1 \sc_dm/sl2/mxl/mux  ( .x(\sc_dm/sl2/mxl/muxout ), .d0(DMEM_d1_i), 
        .sl(n6), .d1(\sc_dm/scn2 ) );
    latn_1 \sc_dm/sl2/mxl/lph1  ( .q(\sc_dm/sl2/l1_q ), .d(
        \sc_dm/sl2/mxl/muxout ), .g(n8) );
    latn_1 \sc_dm/sl1/lph3  ( .q(DMEM_d0_i_sc), .d(\sc_dm/sl1/l1_q ), .g(n3)
         );
    latn_1 \sc_dm/sl1/lph2  ( .q(\sc_dm/scn2 ), .d(\sc_dm/sl1/l1_q ), .g(n15)
         );
    mux2_1 \sc_dm/sl1/mxl/mux  ( .x(\sc_dm/sl1/mxl/muxout ), .d0(DMEM_d0_i), 
        .sl(n7), .d1(\sc_dm/scn1 ) );
    latn_1 \sc_dm/sl1/mxl/lph1  ( .q(\sc_dm/sl1/l1_q ), .d(
        \sc_dm/sl1/mxl/muxout ), .g(n11) );
    latn_1 \sc_dm/sl0/lph3  ( .q(DMEM_eop_i_sc), .d(\sc_dm/sl0/l1_q ), .g(n1)
         );
    latn_1 \sc_dm/sl0/lph2  ( .q(\sc_dm/scn1 ), .d(\sc_dm/sl0/l1_q ), .g(n15)
         );
    mux2_1 \sc_dm/sl0/mxl/mux  ( .x(\sc_dm/sl0/mxl/muxout ), .d0(DMEM_eop_i), 
        .sl(n4), .d1(\scan[1] ) );
    latn_1 \sc_dm/sl0/mxl/lph1  ( .q(\sc_dm/sl0/l1_q ), .d(
        \sc_dm/sl0/mxl/muxout ), .g(n11) );
    latn_1 \sc_im/sl4/lph3  ( .q(IMEM_d3_i_sc), .d(\sc_im/sl4/l1_q ), .g(n1)
         );
    latn_1 \sc_im/sl4/lph2  ( .q(\scan[1] ), .d(\sc_im/sl4/l1_q ), .g(n12) );
    mux2_1 \sc_im/sl4/mxl/mux  ( .x(\sc_im/sl4/mxl/muxout ), .d0(IMEM_d3_i), 
        .sl(n4), .d1(\sc_im/scn4 ) );
    latn_1 \sc_im/sl4/mxl/lph1  ( .q(\sc_im/sl4/l1_q ), .d(
        \sc_im/sl4/mxl/muxout ), .g(n8) );
    latn_1 \sc_im/sl3/lph3  ( .q(IMEM_d2_i_sc), .d(\sc_im/sl3/l1_q ), .g(n1)
         );
    latn_1 \sc_im/sl3/lph2  ( .q(\sc_im/scn4 ), .d(\sc_im/sl3/l1_q ), .g(n14)
         );
    mux2_1 \sc_im/sl3/mxl/mux  ( .x(\sc_im/sl3/mxl/muxout ), .d0(IMEM_d2_i), 
        .sl(n7), .d1(\sc_im/scn3 ) );
    latn_1 \sc_im/sl3/mxl/lph1  ( .q(\sc_im/sl3/l1_q ), .d(
        \sc_im/sl3/mxl/muxout ), .g(n10) );
    latn_1 \sc_im/sl2/lph3  ( .q(IMEM_d1_i_sc), .d(\sc_im/sl2/l1_q ), .g(n1)
         );
    latn_1 \sc_im/sl2/lph2  ( .q(\sc_im/scn3 ), .d(\sc_im/sl2/l1_q ), .g(n14)
         );
    mux2_1 \sc_im/sl2/mxl/mux  ( .x(\sc_im/sl2/mxl/muxout ), .d0(IMEM_d1_i), 
        .sl(n6), .d1(\sc_im/scn2 ) );
    latn_1 \sc_im/sl2/mxl/lph1  ( .q(\sc_im/sl2/l1_q ), .d(
        \sc_im/sl2/mxl/muxout ), .g(n10) );
    latn_1 \sc_im/sl1/lph3  ( .q(IMEM_d0_i_sc), .d(\sc_im/sl1/l1_q ), .g(n1)
         );
    latn_1 \sc_im/sl1/lph2  ( .q(\sc_im/scn2 ), .d(\sc_im/sl1/l1_q ), .g(n12)
         );
    mux2_1 \sc_im/sl1/mxl/mux  ( .x(\sc_im/sl1/mxl/muxout ), .d0(IMEM_d0_i), 
        .sl(n6), .d1(\sc_im/scn1 ) );
    latn_1 \sc_im/sl1/mxl/lph1  ( .q(\sc_im/sl1/l1_q ), .d(
        \sc_im/sl1/mxl/muxout ), .g(n8) );
    latn_1 \sc_im/sl0/lph3  ( .q(IMEM_eop_i_sc), .d(\sc_im/sl0/l1_q ), .g(n1)
         );
    latn_1 \sc_im/sl0/lph2  ( .q(\sc_im/scn1 ), .d(\sc_im/sl0/l1_q ), .g(n14)
         );
    mux2_1 \sc_im/sl0/mxl/mux  ( .x(\sc_im/sl0/mxl/muxout ), .d0(IMEM_eop_i), 
        .sl(n6), .d1(test_si) );
    latn_1 \sc_im/sl0/mxl/lph1  ( .q(\sc_im/sl0/l1_q ), .d(
        \sc_im/sl0/mxl/muxout ), .g(n10) );
    buf_3 U1 ( .x(n5), .a(test_se) );
    buf_1 U2 ( .x(n1), .a(phi3) );
    buf_1 U3 ( .x(n3), .a(phi3) );
    buf_3 U4 ( .x(n2), .a(phi3) );
    buf_3 U5 ( .x(n4), .a(test_se) );
    buf_3 U6 ( .x(n7), .a(test_se) );
    buf_3 U7 ( .x(n6), .a(test_se) );
    buf_3 U8 ( .x(n8), .a(phi1) );
    buf_3 U9 ( .x(n11), .a(phi1) );
    buf_3 U10 ( .x(n9), .a(phi1) );
    buf_3 U11 ( .x(n10), .a(phi1) );
    buf_3 U12 ( .x(n12), .a(phi2) );
    buf_3 U13 ( .x(n15), .a(phi2) );
    buf_3 U14 ( .x(n13), .a(phi2) );
    buf_3 U15 ( .x(n14), .a(phi2) );
endmodule


module wishbone ( reset_b, clk, ch_we_i, ch_dat_i, ch_adr_i, ch_req_i, 
    ch_ack_i, ch_req_o, ch_dat_o, ch_ack_o, wb_we_o, wb_stb_cyc_o, wb_dat_o, 
    wb_adr_o, wb_dat_i, wb_ack_i );
input  [31:0] ch_dat_i;
input  [11:0] ch_adr_i;
output [31:0] ch_dat_o;
output [31:0] wb_dat_o;
output [11:0] wb_adr_o;
input  [31:0] wb_dat_i;
input  reset_b, clk, ch_we_i, ch_req_i, ch_ack_o, wb_ack_i;
output ch_ack_i, ch_req_o, wb_we_o, wb_stb_cyc_o;
    wire \ch_dat_i[31] , \ch_dat_i[30] , \ch_dat_i[29] , \ch_dat_i[28] , 
        \ch_dat_i[27] , \ch_dat_i[26] , \ch_dat_i[25] , \ch_dat_i[24] , 
        \ch_dat_i[23] , \ch_dat_i[22] , \ch_dat_i[21] , \ch_dat_i[20] , 
        \ch_dat_i[19] , \ch_dat_i[18] , \ch_dat_i[17] , \ch_dat_i[16] , 
        \ch_dat_i[15] , \ch_dat_i[14] , \ch_dat_i[13] , \ch_dat_i[12] , 
        \ch_dat_i[11] , \ch_dat_i[10] , \ch_dat_i[9] , \ch_dat_i[8] , 
        \ch_dat_i[7] , \ch_dat_i[6] , \ch_dat_i[5] , \ch_dat_i[4] , 
        \ch_dat_i[3] , \ch_dat_i[2] , \ch_dat_i[1] , \ch_dat_i[0] , 
        \ch_adr_i[11] , \ch_adr_i[10] , \ch_adr_i[9] , \ch_adr_i[8] , 
        \ch_adr_i[7] , \ch_adr_i[6] , \ch_adr_i[5] , \ch_adr_i[4] , 
        \ch_adr_i[3] , \ch_adr_i[2] , \ch_adr_i[1] , \ch_adr_i[0] , 
        ch_req_o_wire, rin1, rsync, sync_ack_l, sync_ack_inv, ch_idle, 
        \reqoGate/nr , \reqoGate/nd , \reqoGate/n2 , n1, n2, n3, n4, n5, n6, 
        n7;
    assign wb_we_o = ch_we_i;
    assign \ch_dat_i[31]  = ch_dat_i[31];
    assign \ch_dat_i[30]  = ch_dat_i[30];
    assign \ch_dat_i[29]  = ch_dat_i[29];
    assign \ch_dat_i[28]  = ch_dat_i[28];
    assign \ch_dat_i[27]  = ch_dat_i[27];
    assign \ch_dat_i[26]  = ch_dat_i[26];
    assign \ch_dat_i[25]  = ch_dat_i[25];
    assign \ch_dat_i[24]  = ch_dat_i[24];
    assign \ch_dat_i[23]  = ch_dat_i[23];
    assign \ch_dat_i[22]  = ch_dat_i[22];
    assign \ch_dat_i[21]  = ch_dat_i[21];
    assign \ch_dat_i[20]  = ch_dat_i[20];
    assign \ch_dat_i[19]  = ch_dat_i[19];
    assign \ch_dat_i[18]  = ch_dat_i[18];
    assign \ch_dat_i[17]  = ch_dat_i[17];
    assign \ch_dat_i[16]  = ch_dat_i[16];
    assign \ch_dat_i[15]  = ch_dat_i[15];
    assign \ch_dat_i[14]  = ch_dat_i[14];
    assign \ch_dat_i[13]  = ch_dat_i[13];
    assign \ch_dat_i[12]  = ch_dat_i[12];
    assign \ch_dat_i[11]  = ch_dat_i[11];
    assign \ch_dat_i[10]  = ch_dat_i[10];
    assign \ch_dat_i[9]  = ch_dat_i[9];
    assign \ch_dat_i[8]  = ch_dat_i[8];
    assign \ch_dat_i[7]  = ch_dat_i[7];
    assign \ch_dat_i[6]  = ch_dat_i[6];
    assign \ch_dat_i[5]  = ch_dat_i[5];
    assign \ch_dat_i[4]  = ch_dat_i[4];
    assign \ch_dat_i[3]  = ch_dat_i[3];
    assign \ch_dat_i[2]  = ch_dat_i[2];
    assign \ch_dat_i[1]  = ch_dat_i[1];
    assign \ch_dat_i[0]  = ch_dat_i[0];
    assign \ch_adr_i[11]  = ch_adr_i[11];
    assign \ch_adr_i[10]  = ch_adr_i[10];
    assign \ch_adr_i[9]  = ch_adr_i[9];
    assign \ch_adr_i[8]  = ch_adr_i[8];
    assign \ch_adr_i[7]  = ch_adr_i[7];
    assign \ch_adr_i[6]  = ch_adr_i[6];
    assign \ch_adr_i[5]  = ch_adr_i[5];
    assign \ch_adr_i[4]  = ch_adr_i[4];
    assign \ch_adr_i[3]  = ch_adr_i[3];
    assign \ch_adr_i[2]  = ch_adr_i[2];
    assign \ch_adr_i[1]  = ch_adr_i[1];
    assign \ch_adr_i[0]  = ch_adr_i[0];
    assign ch_ack_i = ch_req_o;
    assign wb_dat_o[31] = \ch_dat_i[31] ;
    assign wb_dat_o[30] = \ch_dat_i[30] ;
    assign wb_dat_o[29] = \ch_dat_i[29] ;
    assign wb_dat_o[28] = \ch_dat_i[28] ;
    assign wb_dat_o[27] = \ch_dat_i[27] ;
    assign wb_dat_o[26] = \ch_dat_i[26] ;
    assign wb_dat_o[25] = \ch_dat_i[25] ;
    assign wb_dat_o[24] = \ch_dat_i[24] ;
    assign wb_dat_o[23] = \ch_dat_i[23] ;
    assign wb_dat_o[22] = \ch_dat_i[22] ;
    assign wb_dat_o[21] = \ch_dat_i[21] ;
    assign wb_dat_o[20] = \ch_dat_i[20] ;
    assign wb_dat_o[19] = \ch_dat_i[19] ;
    assign wb_dat_o[18] = \ch_dat_i[18] ;
    assign wb_dat_o[17] = \ch_dat_i[17] ;
    assign wb_dat_o[16] = \ch_dat_i[16] ;
    assign wb_dat_o[15] = \ch_dat_i[15] ;
    assign wb_dat_o[14] = \ch_dat_i[14] ;
    assign wb_dat_o[13] = \ch_dat_i[13] ;
    assign wb_dat_o[12] = \ch_dat_i[12] ;
    assign wb_dat_o[11] = \ch_dat_i[11] ;
    assign wb_dat_o[10] = \ch_dat_i[10] ;
    assign wb_dat_o[9] = \ch_dat_i[9] ;
    assign wb_dat_o[8] = \ch_dat_i[8] ;
    assign wb_dat_o[7] = \ch_dat_i[7] ;
    assign wb_dat_o[6] = \ch_dat_i[6] ;
    assign wb_dat_o[5] = \ch_dat_i[5] ;
    assign wb_dat_o[4] = \ch_dat_i[4] ;
    assign wb_dat_o[3] = \ch_dat_i[3] ;
    assign wb_dat_o[2] = \ch_dat_i[2] ;
    assign wb_dat_o[1] = \ch_dat_i[1] ;
    assign wb_dat_o[0] = \ch_dat_i[0] ;
    assign wb_adr_o[11] = \ch_adr_i[11] ;
    assign wb_adr_o[10] = \ch_adr_i[10] ;
    assign wb_adr_o[9] = \ch_adr_i[9] ;
    assign wb_adr_o[8] = \ch_adr_i[8] ;
    assign wb_adr_o[7] = \ch_adr_i[7] ;
    assign wb_adr_o[6] = \ch_adr_i[6] ;
    assign wb_adr_o[5] = \ch_adr_i[5] ;
    assign wb_adr_o[4] = \ch_adr_i[4] ;
    assign wb_adr_o[3] = \ch_adr_i[3] ;
    assign wb_adr_o[2] = \ch_adr_i[2] ;
    assign wb_adr_o[1] = \ch_adr_i[1] ;
    assign wb_adr_o[0] = \ch_adr_i[0] ;
    dffph_2 \ch_dat_o_reg[4]  ( .q(ch_dat_o[4]), .d(wb_dat_i[4]), .ck(n7), .g(
        n4) );
    dffph_2 \ch_dat_o_reg[3]  ( .q(ch_dat_o[3]), .d(wb_dat_i[3]), .ck(n7), .g(
        n4) );
    dffph_2 \ch_dat_o_reg[2]  ( .q(ch_dat_o[2]), .d(wb_dat_i[2]), .ck(n7), .g(
        n4) );
    dffph_2 \ch_dat_o_reg[1]  ( .q(ch_dat_o[1]), .d(wb_dat_i[1]), .ck(n7), .g(
        n4) );
    dffph_2 \ch_dat_o_reg[0]  ( .q(ch_dat_o[0]), .d(wb_dat_i[0]), .ck(n7), .g(
        n3) );
    oa21_2 \reqoGate/U1  ( .x(\reqoGate/n2 ), .a(\reqoGate/n2 ), .b(
        \reqoGate/nr ), .c(\reqoGate/nd ) );
    ao33_1 \cycGate/U1/U1  ( .x(wb_stb_cyc_o), .a(sync_ack_inv), .b(
        wb_stb_cyc_o), .c(reset_b), .d(sync_ack_inv), .e(rsync), .f(ch_idle)
         );
    dffph_2 \ch_dat_o_reg[19]  ( .q(ch_dat_o[19]), .d(wb_dat_i[19]), .ck(n5), 
        .g(n2) );
    dffph_2 \ch_dat_o_reg[18]  ( .q(ch_dat_o[18]), .d(wb_dat_i[18]), .ck(n5), 
        .g(n2) );
    dffph_2 \ch_dat_o_reg[17]  ( .q(ch_dat_o[17]), .d(wb_dat_i[17]), .ck(n6), 
        .g(n2) );
    dffph_2 \ch_dat_o_reg[16]  ( .q(ch_dat_o[16]), .d(wb_dat_i[16]), .ck(n5), 
        .g(n3) );
    dffph_2 \ch_dat_o_reg[15]  ( .q(ch_dat_o[15]), .d(wb_dat_i[15]), .ck(n6), 
        .g(n3) );
    dffph_2 \ch_dat_o_reg[14]  ( .q(ch_dat_o[14]), .d(wb_dat_i[14]), .ck(n6), 
        .g(n3) );
    dffph_2 \ch_dat_o_reg[13]  ( .q(ch_dat_o[13]), .d(wb_dat_i[13]), .ck(n6), 
        .g(n3) );
    dffph_2 \ch_dat_o_reg[12]  ( .q(ch_dat_o[12]), .d(wb_dat_i[12]), .ck(n6), 
        .g(n3) );
    dffph_2 \ch_dat_o_reg[11]  ( .q(ch_dat_o[11]), .d(wb_dat_i[11]), .ck(n7), 
        .g(n4) );
    dffph_2 \ch_dat_o_reg[10]  ( .q(ch_dat_o[10]), .d(wb_dat_i[10]), .ck(n7), 
        .g(n4) );
    dffph_2 \ch_dat_o_reg[9]  ( .q(ch_dat_o[9]), .d(wb_dat_i[9]), .ck(n7), .g(
        n4) );
    dffph_2 \ch_dat_o_reg[8]  ( .q(ch_dat_o[8]), .d(wb_dat_i[8]), .ck(n7), .g(
        n4) );
    dffph_2 \ch_dat_o_reg[7]  ( .q(ch_dat_o[7]), .d(wb_dat_i[7]), .ck(n7), .g(
        n4) );
    dffph_2 \ch_dat_o_reg[6]  ( .q(ch_dat_o[6]), .d(wb_dat_i[6]), .ck(n7), .g(
        n4) );
    dffph_2 \ch_dat_o_reg[5]  ( .q(ch_dat_o[5]), .d(wb_dat_i[5]), .ck(n7), .g(
        n4) );
    dffpr_2 rsync_reg ( .q(rsync), .rb(reset_b), .d(rin1), .ck(n6) );
    dffpr_2 rin1_reg ( .q(rin1), .rb(reset_b), .d(ch_req_i), .ck(n6) );
    dffpr_2 sync_ack_l_reg ( .q(sync_ack_l), .qb(sync_ack_inv), .rb(reset_b), 
        .d(n2), .ck(n6) );
    dffph_2 \ch_dat_o_reg[31]  ( .q(ch_dat_o[31]), .d(wb_dat_i[31]), .ck(n5), 
        .g(n3) );
    dffph_2 \ch_dat_o_reg[30]  ( .q(ch_dat_o[30]), .d(wb_dat_i[30]), .ck(n6), 
        .g(n2) );
    dffph_2 \ch_dat_o_reg[29]  ( .q(ch_dat_o[29]), .d(wb_dat_i[29]), .ck(n5), 
        .g(n3) );
    dffph_2 \ch_dat_o_reg[28]  ( .q(ch_dat_o[28]), .d(wb_dat_i[28]), .ck(n6), 
        .g(n2) );
    dffph_2 \ch_dat_o_reg[27]  ( .q(ch_dat_o[27]), .d(wb_dat_i[27]), .ck(n5), 
        .g(n3) );
    dffph_2 \ch_dat_o_reg[26]  ( .q(ch_dat_o[26]), .d(wb_dat_i[26]), .ck(n6), 
        .g(n2) );
    dffph_2 \ch_dat_o_reg[25]  ( .q(ch_dat_o[25]), .d(wb_dat_i[25]), .ck(n5), 
        .g(n3) );
    dffph_2 \ch_dat_o_reg[24]  ( .q(ch_dat_o[24]), .d(wb_dat_i[24]), .ck(n5), 
        .g(n2) );
    dffph_2 \ch_dat_o_reg[23]  ( .q(ch_dat_o[23]), .d(wb_dat_i[23]), .ck(n5), 
        .g(n3) );
    dffph_2 \ch_dat_o_reg[22]  ( .q(ch_dat_o[22]), .d(wb_dat_i[22]), .ck(n5), 
        .g(n2) );
    dffph_2 \ch_dat_o_reg[21]  ( .q(ch_dat_o[21]), .d(wb_dat_i[21]), .ck(n5), 
        .g(n2) );
    dffph_2 \ch_dat_o_reg[20]  ( .q(ch_dat_o[20]), .d(wb_dat_i[20]), .ck(n5), 
        .g(n2) );
    nor3_0 U3 ( .x(\reqoGate/nr ), .a(n1), .b(sync_ack_l), .c(rsync) );
    nand3_0 U4 ( .x(\reqoGate/nd ), .a(rsync), .b(n1), .c(sync_ack_l) );
    inv_0 U5 ( .x(ch_req_o_wire), .a(\reqoGate/n2 ) );
    nor2_0 U6 ( .x(ch_idle), .a(ch_req_o), .b(ch_ack_o) );
    nor2i_0 U7 ( .x(n1), .a(reset_b), .b(ch_ack_o) );
    buf_3 U8 ( .x(n2), .a(wb_ack_i) );
    buf_3 U9 ( .x(n4), .a(wb_ack_i) );
    buf_3 U10 ( .x(n3), .a(wb_ack_i) );
    buf_3 U11 ( .x(n5), .a(clk) );
    buf_3 U12 ( .x(n7), .a(clk) );
    buf_3 U13 ( .x(n6), .a(clk) );
    buf_3 U14 ( .x(ch_req_o), .a(ch_req_o_wire) );
endmodule


module t_adec_wb ( e_h, e_l, r_h, r_l, e_dp, e_ip, e_tic, r_dp, r_ip, r_tic, 
    tag_h, tag_l );
output [2:0] e_h;
output [2:0] e_l;
output [2:0] r_h;
output [2:0] r_l;
input  [2:0] e_dp;
input  [2:0] e_ip;
input  [2:0] e_tic;
input  [2:0] r_dp;
input  [2:0] r_ip;
input  [2:0] r_tic;
input  [4:0] tag_h;
input  [4:0] tag_l;
    wire \e_l[2] , \e_l[1] , \tag_h[4] , \e_l[0] ;
    assign e_h[2] = 1'b0;
    assign e_h[1] = \e_l[0] ;
    assign e_h[0] = \e_l[1] ;
    assign e_l[2] = \e_l[2] ;
    assign e_l[1] = \e_l[1] ;
    assign e_l[0] = \e_l[0] ;
    assign r_h[2] = \e_l[1] ;
    assign r_h[1] = \tag_h[4] ;
    assign r_h[0] = 1'b0;
    assign r_l[2] = \e_l[0] ;
    assign r_l[0] = \e_l[2] ;
    assign \tag_h[4]  = tag_h[4];
    or2_1 U3 ( .x(r_l[1]), .a(\e_l[0] ), .b(tag_h[3]) );
    buf_3 U6 ( .x(\e_l[0] ), .a(tag_h[2]) );
    or2_2 U7 ( .x(\e_l[2] ), .a(\tag_h[4] ), .b(r_l[1]) );
    or2_2 U8 ( .x(\e_l[1] ), .a(tag_h[3]), .b(\tag_h[4] ) );
endmodule


module chain_sendmux8_4 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/naa , \U1693/bdone , \U1693/net3 , 
        \U1693/drivemonitor , \U1693/net2 , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendmux8_5 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/naa , \U1693/bdone , \U1693/net3 , 
        \U1693/drivemonitor , \U1693/net2 , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendmux8_6 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/naa , \U1693/bdone , \U1693/net3 , 
        \U1693/drivemonitor , \U1693/net2 , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendmux8_7 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/naa , \U1693/bdone , \U1693/net3 , 
        \U1693/drivemonitor , \U1693/net2 , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendword_0 ( ctrlack, oh, ol, chainackff, ctrlreq, ih, il );
output [7:0] oh;
output [7:0] ol;
input  [31:0] ih;
input  [31:0] il;
input  chainackff, ctrlreq;
output ctrlack;
    wire \third_oh[7] , \third_oh[6] , \third_oh[5] , \third_oh[4] , 
        \third_oh[3] , \third_oh[2] , \third_oh[1] , \third_oh[0] , 
        \fourth_ol[7] , \fourth_ol[6] , \fourth_ol[5] , \fourth_ol[4] , 
        \fourth_ol[3] , \fourth_ol[2] , \fourth_ol[1] , \fourth_ol[0] , 
        \third_ol[7] , \third_ol[6] , \third_ol[5] , \third_ol[4] , 
        \third_ol[3] , \third_ol[2] , \third_ol[1] , \third_ol[0] , 
        \fourth_oh[7] , \fourth_oh[6] , \fourth_oh[5] , \fourth_oh[4] , 
        \fourth_oh[3] , \fourth_oh[2] , \fourth_oh[1] , \fourth_oh[0] , 
        \second_oh[7] , \second_oh[6] , \second_oh[5] , \second_oh[4] , 
        \second_oh[3] , \second_oh[2] , \second_oh[1] , \second_oh[0] , 
        \second_ol[7] , \second_ol[6] , \second_ol[5] , \second_ol[4] , 
        \second_ol[3] , \second_ol[2] , \second_ol[1] , \second_ol[0] , 
        \first_oh[7] , \first_oh[6] , \first_oh[5] , \first_oh[4] , 
        \first_oh[3] , \first_oh[2] , \first_oh[1] , \first_oh[0] , 
        \first_ol[7] , \first_ol[6] , \first_ol[5] , \first_ol[4] , 
        \first_ol[3] , \first_ol[2] , \first_ol[1] , \first_ol[0] , net44, 
        net51, net58, bctrlreq, \U309_0_/n5 , \U309_0_/n1 , \U309_0_/n2 , 
        \U309_0_/n3 , \U309_0_/n4 , \U309_1_/n5 , \U309_1_/n1 , \U309_1_/n2 , 
        \U309_1_/n3 , \U309_1_/n4 , \U309_2_/n5 , \U309_2_/n1 , \U309_2_/n2 , 
        \U309_2_/n3 , \U309_2_/n4 , \U309_3_/n5 , \U309_3_/n1 , \U309_3_/n2 , 
        \U309_3_/n3 , \U309_3_/n4 , \U309_4_/n5 , \U309_4_/n1 , \U309_4_/n2 , 
        \U309_4_/n3 , \U309_4_/n4 , \U309_5_/n5 , \U309_5_/n1 , \U309_5_/n2 , 
        \U309_5_/n3 , \U309_5_/n4 , \U309_6_/n5 , \U309_6_/n1 , \U309_6_/n2 , 
        \U309_6_/n3 , \U309_6_/n4 , \U309_7_/n5 , \U309_7_/n1 , \U309_7_/n2 , 
        \U309_7_/n3 , \U309_7_/n4 , \U310_0_/n5 , \U310_0_/n1 , \U310_0_/n2 , 
        \U310_0_/n3 , \U310_0_/n4 , \U310_1_/n5 , \U310_1_/n1 , \U310_1_/n2 , 
        \U310_1_/n3 , \U310_1_/n4 , \U310_2_/n5 , \U310_2_/n1 , \U310_2_/n2 , 
        \U310_2_/n3 , \U310_2_/n4 , \U310_3_/n5 , \U310_3_/n1 , \U310_3_/n2 , 
        \U310_3_/n3 , \U310_3_/n4 , \U310_4_/n5 , \U310_4_/n1 , \U310_4_/n2 , 
        \U310_4_/n3 , \U310_4_/n4 , \U310_5_/n5 , \U310_5_/n1 , \U310_5_/n2 , 
        \U310_5_/n3 , \U310_5_/n4 , \U310_6_/n5 , \U310_6_/n1 , \U310_6_/n2 , 
        \U310_6_/n3 , \U310_6_/n4 , \U310_7_/n5 , \U310_7_/n1 , \U310_7_/n2 , 
        \U310_7_/n3 , \U310_7_/n4 ;
    chain_sendmux8_6 I4 ( .ctrlack(ctrlack), .oh({\fourth_oh[7] , 
        \fourth_oh[6] , \fourth_oh[5] , \fourth_oh[4] , \fourth_oh[3] , 
        \fourth_oh[2] , \fourth_oh[1] , \fourth_oh[0] }), .ol({\fourth_ol[7] , 
        \fourth_ol[6] , \fourth_ol[5] , \fourth_ol[4] , \fourth_ol[3] , 
        \fourth_ol[2] , \fourth_ol[1] , \fourth_ol[0] }), .i_h(ih[7:0]), .i_l(
        il[7:0]), .ctrlreq(net44), .oa(chainackff) );
    chain_sendmux8_5 I3 ( .ctrlack(net44), .oh({\third_oh[7] , \third_oh[6] , 
        \third_oh[5] , \third_oh[4] , \third_oh[3] , \third_oh[2] , 
        \third_oh[1] , \third_oh[0] }), .ol({\third_ol[7] , \third_ol[6] , 
        \third_ol[5] , \third_ol[4] , \third_ol[3] , \third_ol[2] , 
        \third_ol[1] , \third_ol[0] }), .i_h(ih[15:8]), .i_l(il[15:8]), 
        .ctrlreq(net51), .oa(chainackff) );
    chain_sendmux8_4 I2 ( .ctrlack(net51), .oh({\second_oh[7] , \second_oh[6] , 
        \second_oh[5] , \second_oh[4] , \second_oh[3] , \second_oh[2] , 
        \second_oh[1] , \second_oh[0] }), .ol({\second_ol[7] , \second_ol[6] , 
        \second_ol[5] , \second_ol[4] , \second_ol[3] , \second_ol[2] , 
        \second_ol[1] , \second_ol[0] }), .i_h(ih[23:16]), .i_l(il[23:16]), 
        .ctrlreq(net58), .oa(chainackff) );
    chain_sendmux8_7 U320 ( .ctrlack(net58), .oh({\first_oh[7] , \first_oh[6] , 
        \first_oh[5] , \first_oh[4] , \first_oh[3] , \first_oh[2] , 
        \first_oh[1] , \first_oh[0] }), .ol({\first_ol[7] , \first_ol[6] , 
        \first_ol[5] , \first_ol[4] , \first_ol[3] , \first_ol[2] , 
        \first_ol[1] , \first_ol[0] }), .i_h(ih[31:24]), .i_l(il[31:24]), 
        .ctrlreq(bctrlreq), .oa(chainackff) );
    buf_2 \U328/U7  ( .x(bctrlreq), .a(ctrlreq) );
    and4_2 \U309_0_/U24  ( .x(\U309_0_/n5 ), .a(\U309_0_/n1 ), .b(\U309_0_/n2 
        ), .c(\U309_0_/n3 ), .d(\U309_0_/n4 ) );
    inv_1 \U309_0_/U1  ( .x(\U309_0_/n1 ), .a(\fourth_oh[0] ) );
    inv_1 \U309_0_/U2  ( .x(\U309_0_/n2 ), .a(\third_oh[0] ) );
    inv_1 \U309_0_/U3  ( .x(\U309_0_/n3 ), .a(\second_oh[0] ) );
    inv_1 \U309_0_/U4  ( .x(\U309_0_/n4 ), .a(\first_oh[0] ) );
    inv_4 \U309_0_/U5  ( .x(oh[0]), .a(\U309_0_/n5 ) );
    and4_2 \U309_1_/U24  ( .x(\U309_1_/n5 ), .a(\U309_1_/n1 ), .b(\U309_1_/n2 
        ), .c(\U309_1_/n3 ), .d(\U309_1_/n4 ) );
    inv_1 \U309_1_/U1  ( .x(\U309_1_/n1 ), .a(\fourth_oh[1] ) );
    inv_1 \U309_1_/U2  ( .x(\U309_1_/n2 ), .a(\third_oh[1] ) );
    inv_1 \U309_1_/U3  ( .x(\U309_1_/n3 ), .a(\second_oh[1] ) );
    inv_1 \U309_1_/U4  ( .x(\U309_1_/n4 ), .a(\first_oh[1] ) );
    inv_4 \U309_1_/U5  ( .x(oh[1]), .a(\U309_1_/n5 ) );
    and4_2 \U309_2_/U24  ( .x(\U309_2_/n5 ), .a(\U309_2_/n1 ), .b(\U309_2_/n2 
        ), .c(\U309_2_/n3 ), .d(\U309_2_/n4 ) );
    inv_1 \U309_2_/U1  ( .x(\U309_2_/n1 ), .a(\fourth_oh[2] ) );
    inv_1 \U309_2_/U2  ( .x(\U309_2_/n2 ), .a(\third_oh[2] ) );
    inv_1 \U309_2_/U3  ( .x(\U309_2_/n3 ), .a(\second_oh[2] ) );
    inv_1 \U309_2_/U4  ( .x(\U309_2_/n4 ), .a(\first_oh[2] ) );
    inv_4 \U309_2_/U5  ( .x(oh[2]), .a(\U309_2_/n5 ) );
    and4_2 \U309_3_/U24  ( .x(\U309_3_/n5 ), .a(\U309_3_/n1 ), .b(\U309_3_/n2 
        ), .c(\U309_3_/n3 ), .d(\U309_3_/n4 ) );
    inv_1 \U309_3_/U1  ( .x(\U309_3_/n1 ), .a(\fourth_oh[3] ) );
    inv_1 \U309_3_/U2  ( .x(\U309_3_/n2 ), .a(\third_oh[3] ) );
    inv_1 \U309_3_/U3  ( .x(\U309_3_/n3 ), .a(\second_oh[3] ) );
    inv_1 \U309_3_/U4  ( .x(\U309_3_/n4 ), .a(\first_oh[3] ) );
    inv_4 \U309_3_/U5  ( .x(oh[3]), .a(\U309_3_/n5 ) );
    and4_2 \U309_4_/U24  ( .x(\U309_4_/n5 ), .a(\U309_4_/n1 ), .b(\U309_4_/n2 
        ), .c(\U309_4_/n3 ), .d(\U309_4_/n4 ) );
    inv_1 \U309_4_/U1  ( .x(\U309_4_/n1 ), .a(\fourth_oh[4] ) );
    inv_1 \U309_4_/U2  ( .x(\U309_4_/n2 ), .a(\third_oh[4] ) );
    inv_1 \U309_4_/U3  ( .x(\U309_4_/n3 ), .a(\second_oh[4] ) );
    inv_1 \U309_4_/U4  ( .x(\U309_4_/n4 ), .a(\first_oh[4] ) );
    inv_4 \U309_4_/U5  ( .x(oh[4]), .a(\U309_4_/n5 ) );
    and4_2 \U309_5_/U24  ( .x(\U309_5_/n5 ), .a(\U309_5_/n1 ), .b(\U309_5_/n2 
        ), .c(\U309_5_/n3 ), .d(\U309_5_/n4 ) );
    inv_1 \U309_5_/U1  ( .x(\U309_5_/n1 ), .a(\fourth_oh[5] ) );
    inv_1 \U309_5_/U2  ( .x(\U309_5_/n2 ), .a(\third_oh[5] ) );
    inv_1 \U309_5_/U3  ( .x(\U309_5_/n3 ), .a(\second_oh[5] ) );
    inv_1 \U309_5_/U4  ( .x(\U309_5_/n4 ), .a(\first_oh[5] ) );
    inv_4 \U309_5_/U5  ( .x(oh[5]), .a(\U309_5_/n5 ) );
    and4_2 \U309_6_/U24  ( .x(\U309_6_/n5 ), .a(\U309_6_/n1 ), .b(\U309_6_/n2 
        ), .c(\U309_6_/n3 ), .d(\U309_6_/n4 ) );
    inv_1 \U309_6_/U1  ( .x(\U309_6_/n1 ), .a(\fourth_oh[6] ) );
    inv_1 \U309_6_/U2  ( .x(\U309_6_/n2 ), .a(\third_oh[6] ) );
    inv_1 \U309_6_/U3  ( .x(\U309_6_/n3 ), .a(\second_oh[6] ) );
    inv_1 \U309_6_/U4  ( .x(\U309_6_/n4 ), .a(\first_oh[6] ) );
    inv_4 \U309_6_/U5  ( .x(oh[6]), .a(\U309_6_/n5 ) );
    and4_2 \U309_7_/U24  ( .x(\U309_7_/n5 ), .a(\U309_7_/n1 ), .b(\U309_7_/n2 
        ), .c(\U309_7_/n3 ), .d(\U309_7_/n4 ) );
    inv_1 \U309_7_/U1  ( .x(\U309_7_/n1 ), .a(\fourth_oh[7] ) );
    inv_1 \U309_7_/U2  ( .x(\U309_7_/n2 ), .a(\third_oh[7] ) );
    inv_1 \U309_7_/U3  ( .x(\U309_7_/n3 ), .a(\second_oh[7] ) );
    inv_1 \U309_7_/U4  ( .x(\U309_7_/n4 ), .a(\first_oh[7] ) );
    inv_4 \U309_7_/U5  ( .x(oh[7]), .a(\U309_7_/n5 ) );
    and4_2 \U310_0_/U24  ( .x(\U310_0_/n5 ), .a(\U310_0_/n1 ), .b(\U310_0_/n2 
        ), .c(\U310_0_/n3 ), .d(\U310_0_/n4 ) );
    inv_1 \U310_0_/U1  ( .x(\U310_0_/n1 ), .a(\fourth_ol[0] ) );
    inv_1 \U310_0_/U2  ( .x(\U310_0_/n2 ), .a(\third_ol[0] ) );
    inv_1 \U310_0_/U3  ( .x(\U310_0_/n3 ), .a(\second_ol[0] ) );
    inv_1 \U310_0_/U4  ( .x(\U310_0_/n4 ), .a(\first_ol[0] ) );
    inv_4 \U310_0_/U5  ( .x(ol[0]), .a(\U310_0_/n5 ) );
    and4_2 \U310_1_/U24  ( .x(\U310_1_/n5 ), .a(\U310_1_/n1 ), .b(\U310_1_/n2 
        ), .c(\U310_1_/n3 ), .d(\U310_1_/n4 ) );
    inv_1 \U310_1_/U1  ( .x(\U310_1_/n1 ), .a(\fourth_ol[1] ) );
    inv_1 \U310_1_/U2  ( .x(\U310_1_/n2 ), .a(\third_ol[1] ) );
    inv_1 \U310_1_/U3  ( .x(\U310_1_/n3 ), .a(\second_ol[1] ) );
    inv_1 \U310_1_/U4  ( .x(\U310_1_/n4 ), .a(\first_ol[1] ) );
    inv_4 \U310_1_/U5  ( .x(ol[1]), .a(\U310_1_/n5 ) );
    and4_2 \U310_2_/U24  ( .x(\U310_2_/n5 ), .a(\U310_2_/n1 ), .b(\U310_2_/n2 
        ), .c(\U310_2_/n3 ), .d(\U310_2_/n4 ) );
    inv_1 \U310_2_/U1  ( .x(\U310_2_/n1 ), .a(\fourth_ol[2] ) );
    inv_1 \U310_2_/U2  ( .x(\U310_2_/n2 ), .a(\third_ol[2] ) );
    inv_1 \U310_2_/U3  ( .x(\U310_2_/n3 ), .a(\second_ol[2] ) );
    inv_1 \U310_2_/U4  ( .x(\U310_2_/n4 ), .a(\first_ol[2] ) );
    inv_4 \U310_2_/U5  ( .x(ol[2]), .a(\U310_2_/n5 ) );
    and4_2 \U310_3_/U24  ( .x(\U310_3_/n5 ), .a(\U310_3_/n1 ), .b(\U310_3_/n2 
        ), .c(\U310_3_/n3 ), .d(\U310_3_/n4 ) );
    inv_1 \U310_3_/U1  ( .x(\U310_3_/n1 ), .a(\fourth_ol[3] ) );
    inv_1 \U310_3_/U2  ( .x(\U310_3_/n2 ), .a(\third_ol[3] ) );
    inv_1 \U310_3_/U3  ( .x(\U310_3_/n3 ), .a(\second_ol[3] ) );
    inv_1 \U310_3_/U4  ( .x(\U310_3_/n4 ), .a(\first_ol[3] ) );
    inv_4 \U310_3_/U5  ( .x(ol[3]), .a(\U310_3_/n5 ) );
    and4_2 \U310_4_/U24  ( .x(\U310_4_/n5 ), .a(\U310_4_/n1 ), .b(\U310_4_/n2 
        ), .c(\U310_4_/n3 ), .d(\U310_4_/n4 ) );
    inv_1 \U310_4_/U1  ( .x(\U310_4_/n1 ), .a(\fourth_ol[4] ) );
    inv_1 \U310_4_/U2  ( .x(\U310_4_/n2 ), .a(\third_ol[4] ) );
    inv_1 \U310_4_/U3  ( .x(\U310_4_/n3 ), .a(\second_ol[4] ) );
    inv_1 \U310_4_/U4  ( .x(\U310_4_/n4 ), .a(\first_ol[4] ) );
    inv_4 \U310_4_/U5  ( .x(ol[4]), .a(\U310_4_/n5 ) );
    and4_2 \U310_5_/U24  ( .x(\U310_5_/n5 ), .a(\U310_5_/n1 ), .b(\U310_5_/n2 
        ), .c(\U310_5_/n3 ), .d(\U310_5_/n4 ) );
    inv_1 \U310_5_/U1  ( .x(\U310_5_/n1 ), .a(\fourth_ol[5] ) );
    inv_1 \U310_5_/U2  ( .x(\U310_5_/n2 ), .a(\third_ol[5] ) );
    inv_1 \U310_5_/U3  ( .x(\U310_5_/n3 ), .a(\second_ol[5] ) );
    inv_1 \U310_5_/U4  ( .x(\U310_5_/n4 ), .a(\first_ol[5] ) );
    inv_4 \U310_5_/U5  ( .x(ol[5]), .a(\U310_5_/n5 ) );
    and4_2 \U310_6_/U24  ( .x(\U310_6_/n5 ), .a(\U310_6_/n1 ), .b(\U310_6_/n2 
        ), .c(\U310_6_/n3 ), .d(\U310_6_/n4 ) );
    inv_1 \U310_6_/U1  ( .x(\U310_6_/n1 ), .a(\fourth_ol[6] ) );
    inv_1 \U310_6_/U2  ( .x(\U310_6_/n2 ), .a(\third_ol[6] ) );
    inv_1 \U310_6_/U3  ( .x(\U310_6_/n3 ), .a(\second_ol[6] ) );
    inv_1 \U310_6_/U4  ( .x(\U310_6_/n4 ), .a(\first_ol[6] ) );
    inv_4 \U310_6_/U5  ( .x(ol[6]), .a(\U310_6_/n5 ) );
    and4_2 \U310_7_/U24  ( .x(\U310_7_/n5 ), .a(\U310_7_/n1 ), .b(\U310_7_/n2 
        ), .c(\U310_7_/n3 ), .d(\U310_7_/n4 ) );
    inv_1 \U310_7_/U1  ( .x(\U310_7_/n1 ), .a(\fourth_ol[7] ) );
    inv_1 \U310_7_/U2  ( .x(\U310_7_/n2 ), .a(\third_ol[7] ) );
    inv_1 \U310_7_/U3  ( .x(\U310_7_/n3 ), .a(\second_ol[7] ) );
    inv_1 \U310_7_/U4  ( .x(\U310_7_/n4 ), .a(\first_ol[7] ) );
    inv_4 \U310_7_/U5  ( .x(ol[7]), .a(\U310_7_/n5 ) );
endmodule


module chain_selement_ga_63 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_trhdr_0 ( chainff_ack, chainh, chainl, eop, hdrack, normal_ack, 
    notify_ack, read_req, routereq, chain_ff_h, chainack, chainff_l, eopack, 
    err, nReset, normal_response, notify_accept, notify_defer, rcol_h, rcol_l, 
    read_ack, rnw_h, rnw_l, routeack, rsize_h, rsize_l, rtag_h, rtag_l );
output [7:0] chainh;
output [7:0] chainl;
input  [7:0] chain_ff_h;
input  [7:0] chainff_l;
input  [1:0] err;
input  [2:0] rcol_h;
input  [2:0] rcol_l;
input  [1:0] rsize_h;
input  [1:0] rsize_l;
input  [4:0] rtag_h;
input  [4:0] rtag_l;
input  chainack, eopack, nReset, normal_response, notify_accept, notify_defer, 
    read_ack, rnw_h, rnw_l, routeack;
output chainff_ack, eop, hdrack, normal_ack, notify_ack, read_req, routereq;
    wire \net334[0] , \net334[1] , \net334[2] , \net334[4] , \net334[6] , 
        \net334[7] , \net413[0] , \net413[1] , \net413[2] , \net413[3] , 
        \net413[4] , \net413[5] , \net413[6] , \net413[7] , \net413[8] , 
        \net413[9] , \net413[10] , \net413[11] , \net413[12] , \net413[13] , 
        \net413[14] , \net413[15] , \net284[0] , \net284[1] , \net284[2] , 
        \net284[3] , \net284[4] , \net284[5] , \net284[6] , \net284[7] , 
        \net288[0] , \net288[1] , \net288[2] , \net288[3] , \net288[4] , 
        \net288[5] , \net288[6] , \net288[7] , \net343[0] , \net343[1] , 
        \net343[2] , \net343[3] , \net343[5] , \net343[6] , \net343[7] , 
        \hdr[17] , \hdr[16] , \hdr[1] , \hdr[0] , \drive_h[1] , \drive_h[0] , 
        \drive_l[1] , \drive_l[0] , done_write, dowrite, done_eop, ctrl_cd, 
        done_read, done_hdr, done_defer, net321, net362, net359, done_accept, 
        net332, net337, net340, done_pl, net364, donotify, net383, net0230, 
        net407, \U319/U21/U1/loop , \U323/U21/U1/loop , \U320/U21/U1/loop , 
        \U321/U21/U1/loop , \U322/U21/U1/loop , \U311/U28/Z , \U311/U32/Z , 
        \U311/U20/Z , \U311/U29/Z , \U311/U25/Z , \U311/U33/Z , \U311/U21/Z , 
        \U311/U26/Z , \U311/U34/Z , \U311/U30/Z , \U311/U19/Z , \U311/U27/Z , 
        \U311/U35/Z , \U311/U31/Z , \U311/nz[0] , \U311/nz[1] , \U311/x[1] , 
        \U311/y[3] , \U311/y[2] , \U311/x[7] , \U311/x[6] , \U311/x[4] , 
        \U311/y[1] , \U311/x[3] , \U311/x[2] , \U311/y[0] , \U311/x[5] , 
        \U311/x[0] , \U151/Z , \U210/naa , \U210/bdone , \U210/net3 , 
        \U210/drivemonitor , \U210/net2 , \U210/U1702/Z , \I0/naa , \I0/bdone , 
        \I0/net3 , \I0/drivemonitor , \I0/net2 , \I0/U1702/Z ;
    chain_selement_ga_63 U215 ( .Aa(done_eop), .Br(eop), .Ar(done_pl), .Ba(
        eopack) );
    nor2_1 \U308_0_/U5  ( .x(\net413[15] ), .a(\hdr[16] ), .b(\hdr[0] ) );
    nor2_1 \U308_1_/U5  ( .x(\net413[14] ), .a(\hdr[17] ), .b(\hdr[1] ) );
    nor2_1 \U308_2_/U5  ( .x(\net413[13] ), .a(1'b0), .b(routereq) );
    nor2_1 \U308_3_/U5  ( .x(\net413[12] ), .a(routereq), .b(1'b0) );
    nor2_1 \U308_4_/U5  ( .x(\net413[11] ), .a(1'b0), .b(routereq) );
    nor2_1 \U308_5_/U5  ( .x(\net413[10] ), .a(rnw_h), .b(rnw_l) );
    nor2_1 \U308_6_/U5  ( .x(\net413[9] ), .a(rsize_h[0]), .b(rsize_l[0]) );
    nor2_1 \U308_7_/U5  ( .x(\net413[8] ), .a(rsize_h[1]), .b(rsize_l[1]) );
    nor2_1 \U308_8_/U5  ( .x(\net413[7] ), .a(rtag_h[0]), .b(rtag_l[0]) );
    nor2_1 \U308_9_/U5  ( .x(\net413[6] ), .a(rtag_h[1]), .b(rtag_l[1]) );
    nor2_1 \U308_10_/U5  ( .x(\net413[5] ), .a(rtag_h[2]), .b(rtag_l[2]) );
    nor2_1 \U308_11_/U5  ( .x(\net413[4] ), .a(rtag_h[3]), .b(rtag_l[3]) );
    nor2_1 \U308_12_/U5  ( .x(\net413[3] ), .a(rtag_h[4]), .b(rtag_l[4]) );
    nor2_1 \U308_13_/U5  ( .x(\net413[2] ), .a(rcol_h[0]), .b(rcol_l[0]) );
    nor2_1 \U308_14_/U5  ( .x(\net413[1] ), .a(rcol_h[1]), .b(rcol_l[1]) );
    nor2_1 \U308_15_/U5  ( .x(\net413[0] ), .a(rcol_h[2]), .b(rcol_l[2]) );
    or3_1 \U257/U12  ( .x(net364), .a(donotify), .b(dowrite), .c(read_ack) );
    or3_1 \U297/U12  ( .x(net383), .a(done_defer), .b(done_write), .c(
        done_read) );
    and2_2 \U237/U8  ( .x(\hdr[1] ), .a(nReset), .b(normal_response) );
    and2_1 \U307_0_/U8  ( .x(\net343[7] ), .a(\drive_l[0] ), .b(\hdr[0] ) );
    and2_1 \U307_1_/U8  ( .x(\net343[6] ), .a(\drive_l[0] ), .b(\hdr[1] ) );
    and2_1 \U307_2_/U8  ( .x(\net343[5] ), .a(\drive_l[0] ), .b(routereq) );
    and2_1 \U307_4_/U8  ( .x(\net343[3] ), .a(\drive_l[0] ), .b(routereq) );
    and2_1 \U307_5_/U8  ( .x(\net343[2] ), .a(\drive_l[0] ), .b(rnw_l) );
    and2_1 \U307_6_/U8  ( .x(\net343[1] ), .a(\drive_l[0] ), .b(rsize_l[0]) );
    and2_1 \U307_7_/U8  ( .x(\net343[0] ), .a(\drive_l[0] ), .b(rsize_l[1]) );
    and2_1 \U235/U8  ( .x(net340), .a(err[1]), .b(nReset) );
    and2_1 \U236/U8  ( .x(net337), .a(nReset), .b(err[0]) );
    and2_1 \U306_0_/U8  ( .x(\net334[7] ), .a(\hdr[16] ), .b(\drive_l[1] ) );
    and2_1 \U306_1_/U8  ( .x(\net334[6] ), .a(\hdr[17] ), .b(\drive_l[1] ) );
    and2_1 \U306_3_/U8  ( .x(\net334[4] ), .a(routereq), .b(\drive_l[1] ) );
    and2_1 \U306_5_/U8  ( .x(\net334[2] ), .a(rnw_h), .b(\drive_l[1] ) );
    and2_1 \U306_6_/U8  ( .x(\net334[1] ), .a(rsize_h[0]), .b(\drive_l[1] ) );
    and2_1 \U306_7_/U8  ( .x(\net334[0] ), .a(rsize_h[1]), .b(\drive_l[1] ) );
    and2_1 \I1_0_/U8  ( .x(\net284[7] ), .a(rtag_h[0]), .b(\drive_h[1] ) );
    and2_1 \I1_1_/U8  ( .x(\net284[6] ), .a(rtag_h[1]), .b(\drive_h[1] ) );
    and2_1 \I1_2_/U8  ( .x(\net284[5] ), .a(rtag_h[2]), .b(\drive_h[1] ) );
    and2_1 \I1_3_/U8  ( .x(\net284[4] ), .a(rtag_h[3]), .b(\drive_h[1] ) );
    and2_1 \I1_4_/U8  ( .x(\net284[3] ), .a(rtag_h[4]), .b(\drive_h[1] ) );
    and2_1 \I1_5_/U8  ( .x(\net284[2] ), .a(rcol_h[0]), .b(\drive_h[1] ) );
    and2_1 \I1_6_/U8  ( .x(\net284[1] ), .a(rcol_h[1]), .b(\drive_h[1] ) );
    and2_1 \I1_7_/U8  ( .x(\net284[0] ), .a(rcol_h[2]), .b(\drive_h[1] ) );
    and2_1 \I2_0_/U8  ( .x(\net288[7] ), .a(\drive_h[0] ), .b(rtag_l[0]) );
    and2_1 \I2_1_/U8  ( .x(\net288[6] ), .a(\drive_h[0] ), .b(rtag_l[1]) );
    and2_1 \I2_2_/U8  ( .x(\net288[5] ), .a(\drive_h[0] ), .b(rtag_l[2]) );
    and2_1 \I2_3_/U8  ( .x(\net288[4] ), .a(\drive_h[0] ), .b(rtag_l[3]) );
    and2_1 \I2_4_/U8  ( .x(\net288[3] ), .a(\drive_h[0] ), .b(rtag_l[4]) );
    and2_1 \I2_5_/U8  ( .x(\net288[2] ), .a(\drive_h[0] ), .b(rcol_l[0]) );
    and2_1 \I2_6_/U8  ( .x(\net288[1] ), .a(\drive_h[0] ), .b(rcol_l[1]) );
    and2_1 \I2_7_/U8  ( .x(\net288[0] ), .a(\drive_h[0] ), .b(rcol_l[2]) );
    inv_1 \U318/U3  ( .x(net332), .a(routereq) );
    or2_4 \U255/U12  ( .x(notify_ack), .a(done_accept), .b(done_defer) );
    or2_4 \U228/U12  ( .x(\hdr[17] ), .a(notify_defer), .b(notify_accept) );
    or2_4 \U204/U12  ( .x(net321), .a(net359), .b(net362) );
    or2_4 \U221/U12  ( .x(\hdr[16] ), .a(net359), .b(notify_defer) );
    or2_4 \U252/U12  ( .x(normal_ack), .a(done_write), .b(done_read) );
    or2_4 \U280/U12  ( .x(\hdr[0] ), .a(net362), .b(notify_accept) );
    or2_4 \U317/U12  ( .x(routereq), .a(\hdr[17] ), .b(net321) );
    or3_4 \U309_0_/U12  ( .x(chainh[0]), .a(\net334[7] ), .b(\net284[7] ), .c(
        chain_ff_h[0]) );
    or3_4 \U309_1_/U12  ( .x(chainh[1]), .a(\net334[6] ), .b(\net284[6] ), .c(
        chain_ff_h[1]) );
    or3_4 \U309_3_/U12  ( .x(chainh[3]), .a(\net334[4] ), .b(\net284[4] ), .c(
        chain_ff_h[3]) );
    or3_4 \U309_5_/U12  ( .x(chainh[5]), .a(\net334[2] ), .b(\net284[2] ), .c(
        chain_ff_h[5]) );
    or3_4 \U309_6_/U12  ( .x(chainh[6]), .a(\net334[1] ), .b(\net284[1] ), .c(
        chain_ff_h[6]) );
    or3_4 \U309_7_/U12  ( .x(chainh[7]), .a(\net334[0] ), .b(\net284[0] ), .c(
        chain_ff_h[7]) );
    or3_4 \U310_0_/U12  ( .x(chainl[0]), .a(\net343[7] ), .b(\net288[7] ), .c(
        chainff_l[0]) );
    or3_4 \U310_1_/U12  ( .x(chainl[1]), .a(\net343[6] ), .b(\net288[6] ), .c(
        chainff_l[1]) );
    or3_4 \U310_2_/U12  ( .x(chainl[2]), .a(\net343[5] ), .b(\net288[5] ), .c(
        chainff_l[2]) );
    or3_4 \U310_4_/U12  ( .x(chainl[4]), .a(\net343[3] ), .b(\net288[3] ), .c(
        chainff_l[4]) );
    or3_4 \U310_5_/U12  ( .x(chainl[5]), .a(\net343[2] ), .b(\net288[2] ), .c(
        chainff_l[5]) );
    or3_4 \U310_6_/U12  ( .x(chainl[6]), .a(\net343[1] ), .b(\net288[1] ), .c(
        chainff_l[6]) );
    or3_4 \U310_7_/U12  ( .x(chainl[7]), .a(\net343[0] ), .b(\net288[0] ), .c(
        chainff_l[7]) );
    ao222_1 \U311/U37/U18/U1/U1  ( .x(ctrl_cd), .a(\U311/nz[0] ), .b(
        \U311/nz[1] ), .c(\U311/nz[0] ), .d(ctrl_cd), .e(\U311/nz[1] ), .f(
        ctrl_cd) );
    aoi222_1 \U311/U28/U30/U1  ( .x(\U311/x[3] ), .a(\net413[8] ), .b(
        \net413[9] ), .c(\net413[8] ), .d(\U311/U28/Z ), .e(\net413[9] ), .f(
        \U311/U28/Z ) );
    inv_1 \U311/U28/U30/Uinv  ( .x(\U311/U28/Z ), .a(\U311/x[3] ) );
    aoi222_1 \U311/U32/U30/U1  ( .x(\U311/x[0] ), .a(\net413[14] ), .b(
        \net413[15] ), .c(\net413[14] ), .d(\U311/U32/Z ), .e(\net413[15] ), 
        .f(\U311/U32/Z ) );
    inv_1 \U311/U32/U30/Uinv  ( .x(\U311/U32/Z ), .a(\U311/x[0] ) );
    aoi222_1 \U311/U20/U30/U1  ( .x(\U311/x[5] ), .a(\net413[4] ), .b(
        \net413[5] ), .c(\net413[4] ), .d(\U311/U20/Z ), .e(\net413[5] ), .f(
        \U311/U20/Z ) );
    inv_1 \U311/U20/U30/Uinv  ( .x(\U311/U20/Z ), .a(\U311/x[5] ) );
    aoi222_1 \U311/U29/U30/U1  ( .x(\U311/x[2] ), .a(\net413[10] ), .b(
        \net413[11] ), .c(\net413[10] ), .d(\U311/U29/Z ), .e(\net413[11] ), 
        .f(\U311/U29/Z ) );
    inv_1 \U311/U29/U30/Uinv  ( .x(\U311/U29/Z ), .a(\U311/x[2] ) );
    aoi222_1 \U311/U25/U30/U1  ( .x(\U311/x[7] ), .a(\net413[0] ), .b(
        \net413[1] ), .c(\net413[0] ), .d(\U311/U25/Z ), .e(\net413[1] ), .f(
        \U311/U25/Z ) );
    inv_1 \U311/U25/U30/Uinv  ( .x(\U311/U25/Z ), .a(\U311/x[7] ) );
    aoi222_1 \U311/U33/U30/U1  ( .x(\U311/y[0] ), .a(\U311/x[1] ), .b(
        \U311/x[0] ), .c(\U311/x[1] ), .d(\U311/U33/Z ), .e(\U311/x[0] ), .f(
        \U311/U33/Z ) );
    inv_1 \U311/U33/U30/Uinv  ( .x(\U311/U33/Z ), .a(\U311/y[0] ) );
    aoi222_1 \U311/U21/U30/U1  ( .x(\U311/y[2] ), .a(\U311/x[5] ), .b(
        \U311/x[4] ), .c(\U311/x[5] ), .d(\U311/U21/Z ), .e(\U311/x[4] ), .f(
        \U311/U21/Z ) );
    inv_1 \U311/U21/U30/Uinv  ( .x(\U311/U21/Z ), .a(\U311/y[2] ) );
    aoi222_1 \U311/U26/U30/U1  ( .x(\U311/x[6] ), .a(\net413[2] ), .b(
        \net413[3] ), .c(\net413[2] ), .d(\U311/U26/Z ), .e(\net413[3] ), .f(
        \U311/U26/Z ) );
    inv_1 \U311/U26/U30/Uinv  ( .x(\U311/U26/Z ), .a(\U311/x[6] ) );
    aoi222_1 \U311/U34/U30/U1  ( .x(\U311/nz[0] ), .a(\U311/y[1] ), .b(
        \U311/y[0] ), .c(\U311/y[1] ), .d(\U311/U34/Z ), .e(\U311/y[0] ), .f(
        \U311/U34/Z ) );
    inv_1 \U311/U34/U30/Uinv  ( .x(\U311/U34/Z ), .a(\U311/nz[0] ) );
    aoi222_1 \U311/U30/U30/U1  ( .x(\U311/y[1] ), .a(\U311/x[3] ), .b(
        \U311/x[2] ), .c(\U311/x[3] ), .d(\U311/U30/Z ), .e(\U311/x[2] ), .f(
        \U311/U30/Z ) );
    inv_1 \U311/U30/U30/Uinv  ( .x(\U311/U30/Z ), .a(\U311/y[1] ) );
    aoi222_1 \U311/U19/U30/U1  ( .x(\U311/x[4] ), .a(\net413[6] ), .b(
        \net413[7] ), .c(\net413[6] ), .d(\U311/U19/Z ), .e(\net413[7] ), .f(
        \U311/U19/Z ) );
    inv_1 \U311/U19/U30/Uinv  ( .x(\U311/U19/Z ), .a(\U311/x[4] ) );
    aoi222_1 \U311/U27/U30/U1  ( .x(\U311/y[3] ), .a(\U311/x[7] ), .b(
        \U311/x[6] ), .c(\U311/x[7] ), .d(\U311/U27/Z ), .e(\U311/x[6] ), .f(
        \U311/U27/Z ) );
    inv_1 \U311/U27/U30/Uinv  ( .x(\U311/U27/Z ), .a(\U311/y[3] ) );
    aoi222_1 \U311/U35/U30/U1  ( .x(\U311/nz[1] ), .a(\U311/y[3] ), .b(
        \U311/y[2] ), .c(\U311/y[3] ), .d(\U311/U35/Z ), .e(\U311/y[2] ), .f(
        \U311/U35/Z ) );
    inv_1 \U311/U35/U30/Uinv  ( .x(\U311/U35/Z ), .a(\U311/nz[1] ) );
    aoi222_1 \U311/U31/U30/U1  ( .x(\U311/x[1] ), .a(\net413[12] ), .b(
        \net413[13] ), .c(\net413[12] ), .d(\U311/U31/Z ), .e(\net413[13] ), 
        .f(\U311/U31/Z ) );
    inv_1 \U311/U31/U30/Uinv  ( .x(\U311/U31/Z ), .a(\U311/x[1] ) );
    aoi21_1 \U151/U30/U1/U1  ( .x(net407), .a(\U151/Z ), .b(chainff_ack), .c(
        net332) );
    inv_1 \U151/U30/U1/U2  ( .x(\U151/Z ), .a(net407) );
    ao222_1 \U324/U18/U1/U1  ( .x(hdrack), .a(ctrl_cd), .b(net383), .c(ctrl_cd
        ), .d(hdrack), .e(net383), .f(hdrack) );
    ao222_1 \U244/U18/U1/U1  ( .x(donotify), .a(done_hdr), .b(\hdr[17] ), .c(
        done_hdr), .d(donotify), .e(\hdr[17] ), .f(donotify) );
    ao222_1 \U260/U18/U1/U1  ( .x(net362), .a(net337), .b(\hdr[1] ), .c(net337
        ), .d(net362), .e(\hdr[1] ), .f(net362) );
    ao222_1 \U296/U18/U1/U1  ( .x(done_accept), .a(done_eop), .b(notify_accept
        ), .c(done_eop), .d(done_accept), .e(notify_accept), .f(done_accept)
         );
    ao222_1 \U261/U18/U1/U1  ( .x(net359), .a(net340), .b(\hdr[1] ), .c(net340
        ), .d(net359), .e(\hdr[1] ), .f(net359) );
    ao222_1 \U316/U18/U1/U1  ( .x(done_pl), .a(net364), .b(routeack), .c(
        net364), .d(done_pl), .e(routeack), .f(done_pl) );
    ao31_1 \U319/U21/U1/aoi  ( .x(\U319/U21/U1/loop ), .a(\hdr[1] ), .b(
        done_hdr), .c(rnw_h), .d(read_req) );
    oa21_1 \U319/U21/U1/outGate  ( .x(read_req), .a(\hdr[1] ), .b(done_hdr), 
        .c(\U319/U21/U1/loop ) );
    ao31_1 \U323/U21/U1/aoi  ( .x(\U323/U21/U1/loop ), .a(done_eop), .b(
        notify_defer), .c(ctrl_cd), .d(done_defer) );
    oa21_1 \U323/U21/U1/outGate  ( .x(done_defer), .a(done_eop), .b(
        notify_defer), .c(\U323/U21/U1/loop ) );
    ao31_1 \U320/U21/U1/aoi  ( .x(\U320/U21/U1/loop ), .a(\hdr[1] ), .b(
        done_hdr), .c(rnw_l), .d(dowrite) );
    oa21_1 \U320/U21/U1/outGate  ( .x(dowrite), .a(\hdr[1] ), .b(done_hdr), 
        .c(\U320/U21/U1/loop ) );
    ao31_1 \U321/U21/U1/aoi  ( .x(\U321/U21/U1/loop ), .a(read_req), .b(
        done_eop), .c(ctrl_cd), .d(done_read) );
    oa21_1 \U321/U21/U1/outGate  ( .x(done_read), .a(read_req), .b(done_eop), 
        .c(\U321/U21/U1/loop ) );
    ao31_1 \U322/U21/U1/aoi  ( .x(\U322/U21/U1/loop ), .a(dowrite), .b(
        done_eop), .c(ctrl_cd), .d(done_write) );
    oa21_1 \U322/U21/U1/outGate  ( .x(done_write), .a(dowrite), .b(done_eop), 
        .c(\U322/U21/U1/loop ) );
    nor2_2 \U210/U1703/U6  ( .x(done_hdr), .a(\U210/drivemonitor ), .b(
        \U210/naa ) );
    inv_2 \U210/U1699/U3  ( .x(\U210/net2 ), .a(\U210/net3 ) );
    and2_4 \U210/U2_0_/U8  ( .x(\drive_l[0] ), .a(net0230), .b(\U210/net2 ) );
    and2_4 \U210/U2_1_/U8  ( .x(\drive_l[1] ), .a(net0230), .b(\U210/net2 ) );
    inv_1 \U210/U1701/U3  ( .x(\U210/naa ), .a(\U210/bdone ) );
    ao222_1 \U210/U13/U18/U1/U1  ( .x(\U210/drivemonitor ), .a(\drive_l[1] ), 
        .b(\drive_l[0] ), .c(\drive_l[1] ), .d(\U210/drivemonitor ), .e(
        \drive_l[0] ), .f(\U210/drivemonitor ) );
    aoi21_1 \U210/U1702/U30/U1/U1  ( .x(\U210/bdone ), .a(\U210/U1702/Z ), .b(
        chainff_ack), .c(\U210/net2 ) );
    inv_1 \U210/U1702/U30/U1/U2  ( .x(\U210/U1702/Z ), .a(\U210/bdone ) );
    ao23_1 \U210/U1693/U21/U1/U1  ( .x(\U210/net3 ), .a(net0230), .b(
        \U210/net3 ), .c(net0230), .d(\U210/drivemonitor ), .e(chainff_ack) );
    nor2_2 \I0/U1703/U6  ( .x(net0230), .a(\I0/drivemonitor ), .b(\I0/naa ) );
    inv_2 \I0/U1699/U3  ( .x(\I0/net2 ), .a(\I0/net3 ) );
    and2_4 \I0/U2_0_/U8  ( .x(\drive_h[0] ), .a(net407), .b(\I0/net2 ) );
    and2_4 \I0/U2_1_/U8  ( .x(\drive_h[1] ), .a(net407), .b(\I0/net2 ) );
    inv_1 \I0/U1701/U3  ( .x(\I0/naa ), .a(\I0/bdone ) );
    ao222_1 \I0/U13/U18/U1/U1  ( .x(\I0/drivemonitor ), .a(\drive_h[1] ), .b(
        \drive_h[0] ), .c(\drive_h[1] ), .d(\I0/drivemonitor ), .e(
        \drive_h[0] ), .f(\I0/drivemonitor ) );
    aoi21_1 \I0/U1702/U30/U1/U1  ( .x(\I0/bdone ), .a(\I0/U1702/Z ), .b(
        chainff_ack), .c(\I0/net2 ) );
    inv_1 \I0/U1702/U30/U1/U2  ( .x(\I0/U1702/Z ), .a(\I0/bdone ) );
    ao23_1 \I0/U1693/U21/U1/U1  ( .x(\I0/net3 ), .a(net407), .b(\I0/net3 ), 
        .c(net407), .d(\I0/drivemonitor ), .e(chainff_ack) );
    buf_3 U1 ( .x(chainff_ack), .a(chainack) );
    or2_1 U2 ( .x(chainh[4]), .a(chain_ff_h[4]), .b(\net284[3] ) );
    or2_1 U3 ( .x(chainh[2]), .a(chain_ff_h[2]), .b(\net284[5] ) );
    or2_1 U4 ( .x(chainl[3]), .a(chainff_l[3]), .b(\net288[4] ) );
endmodule


module chain_tchdr_0 ( addr_req, col_h, col_l, itag_h, itag_l, lock, ncback, 
    neop, pred, pullcd, reset, rnw_h, rnw_l, seq, size_h, size_l, write_req, 
    chwh, chwl, addr_ack, addr_pull, nReset, nack, write_ack, write_pull );
output [2:0] col_h;
output [2:0] col_l;
output [4:0] itag_h;
output [4:0] itag_l;
output [1:0] lock;
output [1:0] pred;
output [1:0] seq;
output [1:0] size_h;
output [1:0] size_l;
input  [7:0] chwh;
input  [7:0] chwl;
input  addr_ack, addr_pull, nReset, nack, write_ack, write_pull;
output addr_req, ncback, neop, pullcd, reset, rnw_h, rnw_l, write_req;
    wire \ncd[7] , \ncd[6] , \ncd[5] , \ncd[4] , \ncd[3] , \ncd[2] , \ncd[1] , 
        \ncd[0] , net88, receive, pullcdwk, read, net83, ack, net94, n9, 
        \U1664/U28/Z , \U1664/U32/Z , \U1664/U29/Z , \U1664/U33/Z , 
        \U1664/U30/Z , \U1664/U31/Z , \U1664/U37/Z , \U473/Z , \U1664/y[0] , 
        \U1664/y[1] , \U1664/x[1] , \U1664/x[3] , \U1664/x[2] , \U1664/x[0] , 
        \hdr_hld/oh[4] , \hdr_hld/oh[3] , \hdr_hld/ol[4] , \hdr_hld/ol[3] , 
        \hdr_hld/net20 , \hdr_hld/net33 , \hdr_hld/net32 , 
        \hdr_hld/low/drivel , \hdr_hld/low/driveh , \hdr_hld/low/localcd , 
        \hdr_hld/low/ncd[7] , \hdr_hld/low/ncd[6] , \hdr_hld/low/ncd[5] , 
        \hdr_hld/low/ncd[4] , \hdr_hld/low/ncd[3] , \hdr_hld/low/ncd[2] , 
        \hdr_hld/low/ncd[1] , \hdr_hld/low/ncd[0] , \hdr_hld/low/ba , 
        \hdr_hld/low/latch , \hdr_hld/low/acb , \hdr_hld/low/ctrlack_internal , 
        \hdr_hld/low/nlocalcd , \hdr_hld/low/U4/U28/U1/clr , 
        \hdr_hld/low/U4/U28/U1/set , \hdr_hld/low/U1/Z , 
        \hdr_hld/low/U1664/y[0] , \hdr_hld/low/U1664/y[1] , 
        \hdr_hld/low/U1664/x[1] , \hdr_hld/low/U1664/x[3] , 
        \hdr_hld/low/U1664/x[2] , \hdr_hld/low/U1664/x[0] , 
        \hdr_hld/low/U1664/U28/Z , \hdr_hld/low/U1664/U32/Z , 
        \hdr_hld/low/U1664/U29/Z , \hdr_hld/low/U1664/U33/Z , 
        \hdr_hld/low/U1664/U30/Z , \hdr_hld/low/U1664/U31/Z , 
        \hdr_hld/low/U1664/U37/Z , \hdr_hld/low/U1669/nr , 
        \hdr_hld/low/U1669/nd , \hdr_hld/low/U1669/n2 , \hdr_hld/high/drivel , 
        \hdr_hld/high/driveh , \hdr_hld/high/localcd , \hdr_hld/high/ncd[7] , 
        \hdr_hld/high/ncd[6] , \hdr_hld/high/ncd[5] , \hdr_hld/high/ncd[4] , 
        \hdr_hld/high/ncd[3] , \hdr_hld/high/ncd[2] , \hdr_hld/high/ncd[1] , 
        \hdr_hld/high/ncd[0] , \hdr_hld/high/ba , \hdr_hld/high/latch , 
        \hdr_hld/high/acb , \hdr_hld/high/ctrlack_internal , 
        \hdr_hld/high/nlocalcd , \hdr_hld/high/U4/U28/U1/clr , 
        \hdr_hld/high/U4/U28/U1/set , \hdr_hld/high/U1/Z , 
        \hdr_hld/high/U1664/y[0] , \hdr_hld/high/U1664/y[1] , 
        \hdr_hld/high/U1664/x[1] , \hdr_hld/high/U1664/x[3] , 
        \hdr_hld/high/U1664/x[2] , \hdr_hld/high/U1664/x[0] , 
        \hdr_hld/high/U1664/U28/Z , \hdr_hld/high/U1664/U32/Z , 
        \hdr_hld/high/U1664/U29/Z , \hdr_hld/high/U1664/U33/Z , 
        \hdr_hld/high/U1664/U30/Z , \hdr_hld/high/U1664/U31/Z , 
        \hdr_hld/high/U1664/U37/Z , \hdr_hld/high/U1669/nr , 
        \hdr_hld/high/U1669/nd , \hdr_hld/high/U1669/n2 , n1, n2, n3, n4, n5, 
        n6, n7;
    buf_1 U262 ( .x(n9), .a(pullcdwk) );
    or3_2 \U1668/U12  ( .x(ncback), .a(net94), .b(addr_pull), .c(write_pull)
         );
    inv_1 \I0/U3  ( .x(net94), .a(net88) );
    nor2_1 \U514_0_/U5  ( .x(\ncd[0] ), .a(chwh[0]), .b(chwl[0]) );
    nor2_1 \U514_1_/U5  ( .x(\ncd[1] ), .a(chwh[1]), .b(chwl[1]) );
    nor2_1 \U514_2_/U5  ( .x(\ncd[2] ), .a(chwh[2]), .b(chwl[2]) );
    nor2_1 \U514_3_/U5  ( .x(\ncd[3] ), .a(chwh[3]), .b(chwl[3]) );
    nor2_1 \U514_4_/U5  ( .x(\ncd[4] ), .a(chwh[4]), .b(chwl[4]) );
    nor2_1 \U514_5_/U5  ( .x(\ncd[5] ), .a(chwh[5]), .b(chwl[5]) );
    nor2_1 \U514_6_/U5  ( .x(\ncd[6] ), .a(chwh[6]), .b(chwl[6]) );
    nor2_1 \U514_7_/U5  ( .x(\ncd[7] ), .a(chwh[7]), .b(chwl[7]) );
    nor2_1 \U1669/U5  ( .x(neop), .a(read), .b(write_ack) );
    nand2_1 \U303/U5  ( .x(ack), .a(nack), .b(nReset) );
    nand2_1 \U1670/U5  ( .x(net83), .a(neop), .b(nReset) );
    ao222_1 \U47/U18/U1/U1  ( .x(read), .a(addr_ack), .b(rnw_h), .c(addr_ack), 
        .d(read), .e(rnw_h), .f(read) );
    ao222_1 \U48/U18/U1/U1  ( .x(write_req), .a(rnw_l), .b(addr_ack), .c(rnw_l
        ), .d(write_req), .e(addr_ack), .f(write_req) );
    aoi222_1 \U1664/U28/U30/U1  ( .x(\U1664/x[3] ), .a(\ncd[7] ), .b(\ncd[6] ), 
        .c(\ncd[7] ), .d(\U1664/U28/Z ), .e(\ncd[6] ), .f(\U1664/U28/Z ) );
    inv_1 \U1664/U28/U30/Uinv  ( .x(\U1664/U28/Z ), .a(\U1664/x[3] ) );
    aoi222_1 \U1664/U32/U30/U1  ( .x(\U1664/x[0] ), .a(\ncd[1] ), .b(\ncd[0] ), 
        .c(\ncd[1] ), .d(\U1664/U32/Z ), .e(\ncd[0] ), .f(\U1664/U32/Z ) );
    inv_1 \U1664/U32/U30/Uinv  ( .x(\U1664/U32/Z ), .a(\U1664/x[0] ) );
    aoi222_1 \U1664/U29/U30/U1  ( .x(\U1664/x[2] ), .a(\ncd[5] ), .b(\ncd[4] ), 
        .c(\ncd[5] ), .d(\U1664/U29/Z ), .e(\ncd[4] ), .f(\U1664/U29/Z ) );
    inv_1 \U1664/U29/U30/Uinv  ( .x(\U1664/U29/Z ), .a(\U1664/x[2] ) );
    aoi222_1 \U1664/U33/U30/U1  ( .x(\U1664/y[0] ), .a(\U1664/x[1] ), .b(
        \U1664/x[0] ), .c(\U1664/x[1] ), .d(\U1664/U33/Z ), .e(\U1664/x[0] ), 
        .f(\U1664/U33/Z ) );
    inv_1 \U1664/U33/U30/Uinv  ( .x(\U1664/U33/Z ), .a(\U1664/y[0] ) );
    aoi222_1 \U1664/U30/U30/U1  ( .x(\U1664/y[1] ), .a(\U1664/x[3] ), .b(
        \U1664/x[2] ), .c(\U1664/x[3] ), .d(\U1664/U30/Z ), .e(\U1664/x[2] ), 
        .f(\U1664/U30/Z ) );
    inv_1 \U1664/U30/U30/Uinv  ( .x(\U1664/U30/Z ), .a(\U1664/y[1] ) );
    aoi222_1 \U1664/U31/U30/U1  ( .x(\U1664/x[1] ), .a(\ncd[3] ), .b(\ncd[2] ), 
        .c(\ncd[3] ), .d(\U1664/U31/Z ), .e(\ncd[2] ), .f(\U1664/U31/Z ) );
    inv_1 \U1664/U31/U30/Uinv  ( .x(\U1664/U31/Z ), .a(\U1664/x[1] ) );
    aoi222_1 \U1664/U37/U30/U1  ( .x(pullcdwk), .a(\U1664/y[0] ), .b(
        \U1664/y[1] ), .c(\U1664/y[0] ), .d(\U1664/U37/Z ), .e(\U1664/y[1] ), 
        .f(\U1664/U37/Z ) );
    inv_1 \U1664/U37/U30/Uinv  ( .x(\U1664/U37/Z ), .a(pullcdwk) );
    aoi222_1 \U473/U30/U1  ( .x(receive), .a(net83), .b(ack), .c(net83), .d(
        \U473/Z ), .e(ack), .f(\U473/Z ) );
    inv_1 \U473/U30/Uinv  ( .x(\U473/Z ), .a(receive) );
    nor2_1 \hdr_hld/U3/U5  ( .x(net88), .a(\hdr_hld/net32 ), .b(
        \hdr_hld/net33 ) );
    buf_2 \hdr_hld/low/U1653  ( .x(\hdr_hld/low/latch ), .a(\hdr_hld/net32 )
         );
    nor2_1 \hdr_hld/low/U264/U5  ( .x(\hdr_hld/low/nlocalcd ), .a(reset), .b(
        \hdr_hld/low/localcd ) );
    nor2_1 \hdr_hld/low/U1659_0_/U5  ( .x(\hdr_hld/low/ncd[0] ), .a(seq[0]), 
        .b(seq[1]) );
    nor2_1 \hdr_hld/low/U1659_1_/U5  ( .x(\hdr_hld/low/ncd[1] ), .a(pred[0]), 
        .b(pred[1]) );
    nor2_1 \hdr_hld/low/U1659_2_/U5  ( .x(\hdr_hld/low/ncd[2] ), .a(lock[0]), 
        .b(lock[1]) );
    nor2_1 \hdr_hld/low/U1659_3_/U5  ( .x(\hdr_hld/low/ncd[3] ), .a(
        \hdr_hld/ol[3] ), .b(\hdr_hld/oh[3] ) );
    nor2_1 \hdr_hld/low/U1659_4_/U5  ( .x(\hdr_hld/low/ncd[4] ), .a(
        \hdr_hld/ol[4] ), .b(\hdr_hld/oh[4] ) );
    nor2_1 \hdr_hld/low/U1659_5_/U5  ( .x(\hdr_hld/low/ncd[5] ), .a(rnw_l), 
        .b(rnw_h) );
    nor2_1 \hdr_hld/low/U1659_6_/U5  ( .x(\hdr_hld/low/ncd[6] ), .a(size_l[0]), 
        .b(size_h[0]) );
    nor2_1 \hdr_hld/low/U1659_7_/U5  ( .x(\hdr_hld/low/ncd[7] ), .a(size_l[1]), 
        .b(size_h[1]) );
    nor2_1 \hdr_hld/low/U3/U5  ( .x(\hdr_hld/low/ctrlack_internal ), .a(
        \hdr_hld/low/acb ), .b(\hdr_hld/low/ba ) );
    buf_2 \hdr_hld/low/U1665/U7  ( .x(\hdr_hld/low/driveh ), .a(
        \hdr_hld/net20 ) );
    buf_2 \hdr_hld/low/U1666/U7  ( .x(\hdr_hld/low/drivel ), .a(
        \hdr_hld/net20 ) );
    ao23_1 \hdr_hld/low/U1658_0_/U21/U1/U1  ( .x(seq[0]), .a(n7), .b(seq[0]), 
        .c(n7), .d(chwl[0]), .e(n5) );
    ao23_1 \hdr_hld/low/U1658_1_/U21/U1/U1  ( .x(pred[0]), .a(
        \hdr_hld/low/drivel ), .b(pred[0]), .c(\hdr_hld/low/drivel ), .d(chwl
        [1]), .e(n5) );
    ao23_1 \hdr_hld/low/U1658_2_/U21/U1/U1  ( .x(lock[0]), .a(n6), .b(lock[0]), 
        .c(n7), .d(chwl[2]), .e(n5) );
    ao23_1 \hdr_hld/low/U1658_3_/U21/U1/U1  ( .x(\hdr_hld/ol[3] ), .a(
        \hdr_hld/low/drivel ), .b(\hdr_hld/ol[3] ), .c(n6), .d(chwl[3]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_4_/U21/U1/U1  ( .x(\hdr_hld/ol[4] ), .a(n7), .b(
        \hdr_hld/ol[4] ), .c(n6), .d(chwl[4]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_5_/U21/U1/U1  ( .x(rnw_l), .a(n7), .b(rnw_l), 
        .c(n7), .d(chwl[5]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_6_/U21/U1/U1  ( .x(size_l[0]), .a(
        \hdr_hld/low/driveh ), .b(size_l[0]), .c(n6), .d(chwl[6]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_7_/U21/U1/U1  ( .x(size_l[1]), .a(
        \hdr_hld/low/driveh ), .b(size_l[1]), .c(n7), .d(chwl[7]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_0_/U21/U1/U1  ( .x(seq[1]), .a(
        \hdr_hld/low/driveh ), .b(seq[1]), .c(n6), .d(chwh[0]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_1_/U21/U1/U1  ( .x(pred[1]), .a(
        \hdr_hld/low/drivel ), .b(pred[1]), .c(\hdr_hld/low/drivel ), .d(chwh
        [1]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_2_/U21/U1/U1  ( .x(lock[1]), .a(n6), .b(lock[1]), 
        .c(\hdr_hld/low/driveh ), .d(chwh[2]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_3_/U21/U1/U1  ( .x(\hdr_hld/oh[3] ), .a(
        \hdr_hld/low/drivel ), .b(\hdr_hld/oh[3] ), .c(\hdr_hld/low/driveh ), 
        .d(chwh[3]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_4_/U21/U1/U1  ( .x(\hdr_hld/oh[4] ), .a(n7), .b(
        \hdr_hld/oh[4] ), .c(\hdr_hld/low/drivel ), .d(chwh[4]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_5_/U21/U1/U1  ( .x(rnw_h), .a(
        \hdr_hld/low/driveh ), .b(rnw_h), .c(\hdr_hld/low/driveh ), .d(chwh[5]
        ), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_6_/U21/U1/U1  ( .x(size_h[0]), .a(n6), .b(size_h
        [0]), .c(\hdr_hld/low/drivel ), .d(chwh[6]), .e(\hdr_hld/low/latch )
         );
    ao23_1 \hdr_hld/low/U1651_7_/U21/U1/U1  ( .x(size_h[1]), .a(n6), .b(size_h
        [1]), .c(\hdr_hld/low/driveh ), .d(chwh[7]), .e(\hdr_hld/low/latch )
         );
    aoai211_1 \hdr_hld/low/U4/U28/U1/U1  ( .x(\hdr_hld/low/U4/U28/U1/clr ), 
        .a(\hdr_hld/net20 ), .b(\hdr_hld/low/acb ), .c(\hdr_hld/low/nlocalcd ), 
        .d(\hdr_hld/net32 ) );
    nand3_1 \hdr_hld/low/U4/U28/U1/U2  ( .x(\hdr_hld/low/U4/U28/U1/set ), .a(
        \hdr_hld/low/nlocalcd ), .b(\hdr_hld/net20 ), .c(\hdr_hld/low/acb ) );
    nand2_2 \hdr_hld/low/U4/U28/U1/U3  ( .x(\hdr_hld/net32 ), .a(
        \hdr_hld/low/U4/U28/U1/clr ), .b(\hdr_hld/low/U4/U28/U1/set ) );
    oai21_1 \hdr_hld/low/U1/U30/U1/U1  ( .x(\hdr_hld/low/acb ), .a(
        \hdr_hld/low/U1/Z ), .b(\hdr_hld/low/ba ), .c(\hdr_hld/net20 ) );
    inv_1 \hdr_hld/low/U1/U30/U1/U2  ( .x(\hdr_hld/low/U1/Z ), .a(
        \hdr_hld/low/acb ) );
    ao222_1 \hdr_hld/low/U5/U18/U1/U1  ( .x(\hdr_hld/low/ba ), .a(
        \hdr_hld/low/latch ), .b(n9), .c(\hdr_hld/low/latch ), .d(
        \hdr_hld/low/ba ), .e(n9), .f(\hdr_hld/low/ba ) );
    aoi222_1 \hdr_hld/low/U1664/U28/U30/U1  ( .x(\hdr_hld/low/U1664/x[3] ), 
        .a(\hdr_hld/low/ncd[7] ), .b(\hdr_hld/low/ncd[6] ), .c(
        \hdr_hld/low/ncd[7] ), .d(\hdr_hld/low/U1664/U28/Z ), .e(
        \hdr_hld/low/ncd[6] ), .f(\hdr_hld/low/U1664/U28/Z ) );
    inv_1 \hdr_hld/low/U1664/U28/U30/Uinv  ( .x(\hdr_hld/low/U1664/U28/Z ), 
        .a(\hdr_hld/low/U1664/x[3] ) );
    aoi222_1 \hdr_hld/low/U1664/U32/U30/U1  ( .x(\hdr_hld/low/U1664/x[0] ), 
        .a(\hdr_hld/low/ncd[1] ), .b(\hdr_hld/low/ncd[0] ), .c(
        \hdr_hld/low/ncd[1] ), .d(\hdr_hld/low/U1664/U32/Z ), .e(
        \hdr_hld/low/ncd[0] ), .f(\hdr_hld/low/U1664/U32/Z ) );
    inv_1 \hdr_hld/low/U1664/U32/U30/Uinv  ( .x(\hdr_hld/low/U1664/U32/Z ), 
        .a(\hdr_hld/low/U1664/x[0] ) );
    aoi222_1 \hdr_hld/low/U1664/U29/U30/U1  ( .x(\hdr_hld/low/U1664/x[2] ), 
        .a(\hdr_hld/low/ncd[5] ), .b(\hdr_hld/low/ncd[4] ), .c(
        \hdr_hld/low/ncd[5] ), .d(\hdr_hld/low/U1664/U29/Z ), .e(
        \hdr_hld/low/ncd[4] ), .f(\hdr_hld/low/U1664/U29/Z ) );
    inv_1 \hdr_hld/low/U1664/U29/U30/Uinv  ( .x(\hdr_hld/low/U1664/U29/Z ), 
        .a(\hdr_hld/low/U1664/x[2] ) );
    aoi222_1 \hdr_hld/low/U1664/U33/U30/U1  ( .x(\hdr_hld/low/U1664/y[0] ), 
        .a(\hdr_hld/low/U1664/x[1] ), .b(\hdr_hld/low/U1664/x[0] ), .c(
        \hdr_hld/low/U1664/x[1] ), .d(\hdr_hld/low/U1664/U33/Z ), .e(
        \hdr_hld/low/U1664/x[0] ), .f(\hdr_hld/low/U1664/U33/Z ) );
    inv_1 \hdr_hld/low/U1664/U33/U30/Uinv  ( .x(\hdr_hld/low/U1664/U33/Z ), 
        .a(\hdr_hld/low/U1664/y[0] ) );
    aoi222_1 \hdr_hld/low/U1664/U30/U30/U1  ( .x(\hdr_hld/low/U1664/y[1] ), 
        .a(\hdr_hld/low/U1664/x[3] ), .b(\hdr_hld/low/U1664/x[2] ), .c(
        \hdr_hld/low/U1664/x[3] ), .d(\hdr_hld/low/U1664/U30/Z ), .e(
        \hdr_hld/low/U1664/x[2] ), .f(\hdr_hld/low/U1664/U30/Z ) );
    inv_1 \hdr_hld/low/U1664/U30/U30/Uinv  ( .x(\hdr_hld/low/U1664/U30/Z ), 
        .a(\hdr_hld/low/U1664/y[1] ) );
    aoi222_1 \hdr_hld/low/U1664/U31/U30/U1  ( .x(\hdr_hld/low/U1664/x[1] ), 
        .a(\hdr_hld/low/ncd[3] ), .b(\hdr_hld/low/ncd[2] ), .c(
        \hdr_hld/low/ncd[3] ), .d(\hdr_hld/low/U1664/U31/Z ), .e(
        \hdr_hld/low/ncd[2] ), .f(\hdr_hld/low/U1664/U31/Z ) );
    inv_1 \hdr_hld/low/U1664/U31/U30/Uinv  ( .x(\hdr_hld/low/U1664/U31/Z ), 
        .a(\hdr_hld/low/U1664/x[1] ) );
    aoi222_1 \hdr_hld/low/U1664/U37/U30/U1  ( .x(\hdr_hld/low/localcd ), .a(
        \hdr_hld/low/U1664/y[0] ), .b(\hdr_hld/low/U1664/y[1] ), .c(
        \hdr_hld/low/U1664/y[0] ), .d(\hdr_hld/low/U1664/U37/Z ), .e(
        \hdr_hld/low/U1664/y[1] ), .f(\hdr_hld/low/U1664/U37/Z ) );
    inv_1 \hdr_hld/low/U1664/U37/U30/Uinv  ( .x(\hdr_hld/low/U1664/U37/Z ), 
        .a(\hdr_hld/low/localcd ) );
    nor3_1 \hdr_hld/low/U1669/Unr  ( .x(\hdr_hld/low/U1669/nr ), .a(
        \hdr_hld/low/ctrlack_internal ), .b(\hdr_hld/low/drivel ), .c(n6) );
    nand3_1 \hdr_hld/low/U1669/Und  ( .x(\hdr_hld/low/U1669/nd ), .a(
        \hdr_hld/low/ctrlack_internal ), .b(n7), .c(\hdr_hld/low/driveh ) );
    oa21_1 \hdr_hld/low/U1669/U1  ( .x(\hdr_hld/low/U1669/n2 ), .a(
        \hdr_hld/low/U1669/n2 ), .b(\hdr_hld/low/U1669/nr ), .c(
        \hdr_hld/low/U1669/nd ) );
    inv_2 \hdr_hld/low/U1669/U3  ( .x(addr_req), .a(\hdr_hld/low/U1669/n2 ) );
    buf_2 \hdr_hld/high/U1653  ( .x(\hdr_hld/high/latch ), .a(\hdr_hld/net33 )
         );
    nor2_1 \hdr_hld/high/U264/U5  ( .x(\hdr_hld/high/nlocalcd ), .a(reset), 
        .b(\hdr_hld/high/localcd ) );
    nor2_1 \hdr_hld/high/U1659_0_/U5  ( .x(\hdr_hld/high/ncd[0] ), .a(itag_l
        [0]), .b(itag_h[0]) );
    nor2_1 \hdr_hld/high/U1659_1_/U5  ( .x(\hdr_hld/high/ncd[1] ), .a(itag_l
        [1]), .b(itag_h[1]) );
    nor2_1 \hdr_hld/high/U1659_2_/U5  ( .x(\hdr_hld/high/ncd[2] ), .a(itag_l
        [2]), .b(itag_h[2]) );
    nor2_1 \hdr_hld/high/U1659_3_/U5  ( .x(\hdr_hld/high/ncd[3] ), .a(itag_l
        [3]), .b(itag_h[3]) );
    nor2_1 \hdr_hld/high/U1659_4_/U5  ( .x(\hdr_hld/high/ncd[4] ), .a(itag_l
        [4]), .b(itag_h[4]) );
    nor2_1 \hdr_hld/high/U1659_5_/U5  ( .x(\hdr_hld/high/ncd[5] ), .a(col_l[0]
        ), .b(col_h[0]) );
    nor2_1 \hdr_hld/high/U1659_6_/U5  ( .x(\hdr_hld/high/ncd[6] ), .a(col_l[1]
        ), .b(col_h[1]) );
    nor2_1 \hdr_hld/high/U1659_7_/U5  ( .x(\hdr_hld/high/ncd[7] ), .a(col_l[2]
        ), .b(col_h[2]) );
    nor2_1 \hdr_hld/high/U3/U5  ( .x(\hdr_hld/high/ctrlack_internal ), .a(
        \hdr_hld/high/acb ), .b(\hdr_hld/high/ba ) );
    buf_2 \hdr_hld/high/U1665/U7  ( .x(\hdr_hld/high/driveh ), .a(receive) );
    buf_2 \hdr_hld/high/U1666/U7  ( .x(\hdr_hld/high/drivel ), .a(receive) );
    ao23_1 \hdr_hld/high/U1658_0_/U21/U1/U1  ( .x(itag_l[0]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[0]), .c(\hdr_hld/high/drivel ), .d(
        chwl[0]), .e(n1) );
    ao23_1 \hdr_hld/high/U1658_1_/U21/U1/U1  ( .x(itag_l[1]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[1]), .c(\hdr_hld/high/drivel ), .d(
        chwl[1]), .e(n1) );
    ao23_1 \hdr_hld/high/U1658_2_/U21/U1/U1  ( .x(itag_l[2]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[2]), .c(\hdr_hld/high/drivel ), .d(
        chwl[2]), .e(n1) );
    ao23_1 \hdr_hld/high/U1658_3_/U21/U1/U1  ( .x(itag_l[3]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[3]), .c(\hdr_hld/high/drivel ), .d(
        chwl[3]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1658_4_/U21/U1/U1  ( .x(itag_l[4]), .a(n4), .b(
        itag_l[4]), .c(\hdr_hld/high/drivel ), .d(chwl[4]), .e(
        \hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1658_5_/U21/U1/U1  ( .x(col_l[0]), .a(n4), .b(col_l
        [0]), .c(\hdr_hld/high/drivel ), .d(chwl[5]), .e(\hdr_hld/high/latch )
         );
    ao23_1 \hdr_hld/high/U1658_6_/U21/U1/U1  ( .x(col_l[1]), .a(
        \hdr_hld/high/drivel ), .b(col_l[1]), .c(\hdr_hld/high/drivel ), .d(
        chwl[6]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1658_7_/U21/U1/U1  ( .x(col_l[2]), .a(n4), .b(col_l
        [2]), .c(\hdr_hld/high/drivel ), .d(chwl[7]), .e(\hdr_hld/high/latch )
         );
    ao23_1 \hdr_hld/high/U1651_0_/U21/U1/U1  ( .x(itag_h[0]), .a(n2), .b(
        itag_h[0]), .c(n2), .d(chwh[0]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_1_/U21/U1/U1  ( .x(itag_h[1]), .a(n2), .b(
        itag_h[1]), .c(n3), .d(chwh[1]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_2_/U21/U1/U1  ( .x(itag_h[2]), .a(n2), .b(
        itag_h[2]), .c(n3), .d(chwh[2]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_3_/U21/U1/U1  ( .x(itag_h[3]), .a(n2), .b(
        itag_h[3]), .c(n3), .d(chwh[3]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_4_/U21/U1/U1  ( .x(itag_h[4]), .a(n2), .b(
        itag_h[4]), .c(n3), .d(chwh[4]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_5_/U21/U1/U1  ( .x(col_h[0]), .a(n2), .b(col_h
        [0]), .c(n3), .d(chwh[5]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_6_/U21/U1/U1  ( .x(col_h[1]), .a(n2), .b(col_h
        [1]), .c(n2), .d(chwh[6]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_7_/U21/U1/U1  ( .x(col_h[2]), .a(n2), .b(col_h
        [2]), .c(n2), .d(chwh[7]), .e(\hdr_hld/high/latch ) );
    aoai211_1 \hdr_hld/high/U4/U28/U1/U1  ( .x(\hdr_hld/high/U4/U28/U1/clr ), 
        .a(receive), .b(\hdr_hld/high/acb ), .c(\hdr_hld/high/nlocalcd ), .d(
        \hdr_hld/net33 ) );
    nand3_1 \hdr_hld/high/U4/U28/U1/U2  ( .x(\hdr_hld/high/U4/U28/U1/set ), 
        .a(\hdr_hld/high/nlocalcd ), .b(receive), .c(\hdr_hld/high/acb ) );
    nand2_2 \hdr_hld/high/U4/U28/U1/U3  ( .x(\hdr_hld/net33 ), .a(
        \hdr_hld/high/U4/U28/U1/clr ), .b(\hdr_hld/high/U4/U28/U1/set ) );
    oai21_1 \hdr_hld/high/U1/U30/U1/U1  ( .x(\hdr_hld/high/acb ), .a(
        \hdr_hld/high/U1/Z ), .b(\hdr_hld/high/ba ), .c(receive) );
    inv_1 \hdr_hld/high/U1/U30/U1/U2  ( .x(\hdr_hld/high/U1/Z ), .a(
        \hdr_hld/high/acb ) );
    ao222_1 \hdr_hld/high/U5/U18/U1/U1  ( .x(\hdr_hld/high/ba ), .a(
        \hdr_hld/high/latch ), .b(n9), .c(\hdr_hld/high/latch ), .d(
        \hdr_hld/high/ba ), .e(n9), .f(\hdr_hld/high/ba ) );
    aoi222_1 \hdr_hld/high/U1664/U28/U30/U1  ( .x(\hdr_hld/high/U1664/x[3] ), 
        .a(\hdr_hld/high/ncd[7] ), .b(\hdr_hld/high/ncd[6] ), .c(
        \hdr_hld/high/ncd[7] ), .d(\hdr_hld/high/U1664/U28/Z ), .e(
        \hdr_hld/high/ncd[6] ), .f(\hdr_hld/high/U1664/U28/Z ) );
    inv_1 \hdr_hld/high/U1664/U28/U30/Uinv  ( .x(\hdr_hld/high/U1664/U28/Z ), 
        .a(\hdr_hld/high/U1664/x[3] ) );
    aoi222_1 \hdr_hld/high/U1664/U32/U30/U1  ( .x(\hdr_hld/high/U1664/x[0] ), 
        .a(\hdr_hld/high/ncd[1] ), .b(\hdr_hld/high/ncd[0] ), .c(
        \hdr_hld/high/ncd[1] ), .d(\hdr_hld/high/U1664/U32/Z ), .e(
        \hdr_hld/high/ncd[0] ), .f(\hdr_hld/high/U1664/U32/Z ) );
    inv_1 \hdr_hld/high/U1664/U32/U30/Uinv  ( .x(\hdr_hld/high/U1664/U32/Z ), 
        .a(\hdr_hld/high/U1664/x[0] ) );
    aoi222_1 \hdr_hld/high/U1664/U29/U30/U1  ( .x(\hdr_hld/high/U1664/x[2] ), 
        .a(\hdr_hld/high/ncd[5] ), .b(\hdr_hld/high/ncd[4] ), .c(
        \hdr_hld/high/ncd[5] ), .d(\hdr_hld/high/U1664/U29/Z ), .e(
        \hdr_hld/high/ncd[4] ), .f(\hdr_hld/high/U1664/U29/Z ) );
    inv_1 \hdr_hld/high/U1664/U29/U30/Uinv  ( .x(\hdr_hld/high/U1664/U29/Z ), 
        .a(\hdr_hld/high/U1664/x[2] ) );
    aoi222_1 \hdr_hld/high/U1664/U33/U30/U1  ( .x(\hdr_hld/high/U1664/y[0] ), 
        .a(\hdr_hld/high/U1664/x[1] ), .b(\hdr_hld/high/U1664/x[0] ), .c(
        \hdr_hld/high/U1664/x[1] ), .d(\hdr_hld/high/U1664/U33/Z ), .e(
        \hdr_hld/high/U1664/x[0] ), .f(\hdr_hld/high/U1664/U33/Z ) );
    inv_1 \hdr_hld/high/U1664/U33/U30/Uinv  ( .x(\hdr_hld/high/U1664/U33/Z ), 
        .a(\hdr_hld/high/U1664/y[0] ) );
    aoi222_1 \hdr_hld/high/U1664/U30/U30/U1  ( .x(\hdr_hld/high/U1664/y[1] ), 
        .a(\hdr_hld/high/U1664/x[3] ), .b(\hdr_hld/high/U1664/x[2] ), .c(
        \hdr_hld/high/U1664/x[3] ), .d(\hdr_hld/high/U1664/U30/Z ), .e(
        \hdr_hld/high/U1664/x[2] ), .f(\hdr_hld/high/U1664/U30/Z ) );
    inv_1 \hdr_hld/high/U1664/U30/U30/Uinv  ( .x(\hdr_hld/high/U1664/U30/Z ), 
        .a(\hdr_hld/high/U1664/y[1] ) );
    aoi222_1 \hdr_hld/high/U1664/U31/U30/U1  ( .x(\hdr_hld/high/U1664/x[1] ), 
        .a(\hdr_hld/high/ncd[3] ), .b(\hdr_hld/high/ncd[2] ), .c(
        \hdr_hld/high/ncd[3] ), .d(\hdr_hld/high/U1664/U31/Z ), .e(
        \hdr_hld/high/ncd[2] ), .f(\hdr_hld/high/U1664/U31/Z ) );
    inv_1 \hdr_hld/high/U1664/U31/U30/Uinv  ( .x(\hdr_hld/high/U1664/U31/Z ), 
        .a(\hdr_hld/high/U1664/x[1] ) );
    aoi222_1 \hdr_hld/high/U1664/U37/U30/U1  ( .x(\hdr_hld/high/localcd ), .a(
        \hdr_hld/high/U1664/y[0] ), .b(\hdr_hld/high/U1664/y[1] ), .c(
        \hdr_hld/high/U1664/y[0] ), .d(\hdr_hld/high/U1664/U37/Z ), .e(
        \hdr_hld/high/U1664/y[1] ), .f(\hdr_hld/high/U1664/U37/Z ) );
    inv_1 \hdr_hld/high/U1664/U37/U30/Uinv  ( .x(\hdr_hld/high/U1664/U37/Z ), 
        .a(\hdr_hld/high/localcd ) );
    nor3_1 \hdr_hld/high/U1669/Unr  ( .x(\hdr_hld/high/U1669/nr ), .a(
        \hdr_hld/high/ctrlack_internal ), .b(\hdr_hld/high/drivel ), .c(n3) );
    nand3_1 \hdr_hld/high/U1669/Und  ( .x(\hdr_hld/high/U1669/nd ), .a(
        \hdr_hld/high/ctrlack_internal ), .b(\hdr_hld/high/drivel ), .c(n3) );
    oa21_1 \hdr_hld/high/U1669/U1  ( .x(\hdr_hld/high/U1669/n2 ), .a(
        \hdr_hld/high/U1669/n2 ), .b(\hdr_hld/high/U1669/nr ), .c(
        \hdr_hld/high/U1669/nd ) );
    inv_2 \hdr_hld/high/U1669/U3  ( .x(\hdr_hld/net20 ), .a(
        \hdr_hld/high/U1669/n2 ) );
    buf_1 U1 ( .x(n1), .a(\hdr_hld/high/latch ) );
    buf_3 U2 ( .x(n2), .a(\hdr_hld/high/driveh ) );
    buf_3 U3 ( .x(n3), .a(\hdr_hld/high/driveh ) );
    buf_1 U4 ( .x(n4), .a(\hdr_hld/high/drivel ) );
    buf_1 U5 ( .x(n5), .a(\hdr_hld/low/latch ) );
    buf_2 U6 ( .x(n7), .a(\hdr_hld/net20 ) );
    buf_2 U7 ( .x(n6), .a(\hdr_hld/net20 ) );
    inv_2 U8 ( .x(reset), .a(nReset) );
    buf_3 U9 ( .x(pullcd), .a(n9) );
endmodule


module chain_irdemux_32new_0 ( ctrlack, oh, ol, pullreq, pull_h, pull_l, 
    pullcd, reset, ctrlreq );
output [31:0] oh;
output [31:0] ol;
input  [7:0] pull_h;
input  [7:0] pull_l;
input  pullcd, reset, ctrlreq;
output ctrlack, pullreq;
    wire net30, net31, net17, \I0/net20 , \I0/net33 , \I0/net32 , 
        \I0/low/drivel , \I0/low/driveh , \I0/low/localcd , \I0/low/ncd[7] , 
        \I0/low/ncd[6] , \I0/low/ncd[5] , \I0/low/ncd[4] , \I0/low/ncd[3] , 
        \I0/low/ncd[2] , \I0/low/ncd[1] , \I0/low/ncd[0] , \I0/low/ba , 
        \I0/low/latch , \I0/low/acb , \I0/low/ctrlack_internal , 
        \I0/low/nlocalcd , \I0/low/U4/U28/U1/clr , \I0/low/U4/U28/U1/set , 
        \I0/low/U1/Z , \I0/low/U1664/y[0] , \I0/low/U1664/y[1] , 
        \I0/low/U1664/x[1] , \I0/low/U1664/x[3] , \I0/low/U1664/x[2] , 
        \I0/low/U1664/x[0] , \I0/low/U1664/U28/Z , \I0/low/U1664/U32/Z , 
        \I0/low/U1664/U29/Z , \I0/low/U1664/U33/Z , \I0/low/U1664/U30/Z , 
        \I0/low/U1664/U31/Z , \I0/low/U1664/U37/Z , \I0/low/U1669/nr , 
        \I0/low/U1669/nd , \I0/low/U1669/n2 , \I0/high/drivel , 
        \I0/high/driveh , \I0/high/localcd , \I0/high/ncd[7] , 
        \I0/high/ncd[6] , \I0/high/ncd[5] , \I0/high/ncd[4] , \I0/high/ncd[3] , 
        \I0/high/ncd[2] , \I0/high/ncd[1] , \I0/high/ncd[0] , \I0/high/ba , 
        \I0/high/latch , \I0/high/acb , \I0/high/ctrlack_internal , 
        \I0/high/nlocalcd , \I0/high/U4/U28/U1/clr , \I0/high/U4/U28/U1/set , 
        \I0/high/U1/Z , \I0/high/U1664/y[0] , \I0/high/U1664/y[1] , 
        \I0/high/U1664/x[1] , \I0/high/U1664/x[3] , \I0/high/U1664/x[2] , 
        \I0/high/U1664/x[0] , \I0/high/U1664/U28/Z , \I0/high/U1664/U32/Z , 
        \I0/high/U1664/U29/Z , \I0/high/U1664/U33/Z , \I0/high/U1664/U30/Z , 
        \I0/high/U1664/U31/Z , \I0/high/U1664/U37/Z , \I0/high/U1669/nr , 
        \I0/high/U1669/nd , \I0/high/U1669/n2 , \I1/net20 , \I1/net33 , 
        \I1/net32 , \I1/low/drivel , \I1/low/driveh , \I1/low/localcd , 
        \I1/low/ncd[7] , \I1/low/ncd[6] , \I1/low/ncd[5] , \I1/low/ncd[4] , 
        \I1/low/ncd[3] , \I1/low/ncd[2] , \I1/low/ncd[1] , \I1/low/ncd[0] , 
        \I1/low/ba , \I1/low/latch , \I1/low/acb , \I1/low/ctrlack_internal , 
        \I1/low/nlocalcd , \I1/low/U4/U28/U1/clr , \I1/low/U4/U28/U1/set , 
        \I1/low/U1/Z , \I1/low/U1664/y[0] , \I1/low/U1664/y[1] , 
        \I1/low/U1664/x[1] , \I1/low/U1664/x[3] , \I1/low/U1664/x[2] , 
        \I1/low/U1664/x[0] , \I1/low/U1664/U28/Z , \I1/low/U1664/U32/Z , 
        \I1/low/U1664/U29/Z , \I1/low/U1664/U33/Z , \I1/low/U1664/U30/Z , 
        \I1/low/U1664/U31/Z , \I1/low/U1664/U37/Z , \I1/low/U1669/nr , 
        \I1/low/U1669/nd , \I1/low/U1669/n2 , \I1/high/drivel , 
        \I1/high/driveh , \I1/high/localcd , \I1/high/ncd[7] , 
        \I1/high/ncd[6] , \I1/high/ncd[5] , \I1/high/ncd[4] , \I1/high/ncd[3] , 
        \I1/high/ncd[2] , \I1/high/ncd[1] , \I1/high/ncd[0] , \I1/high/ba , 
        \I1/high/latch , \I1/high/acb , \I1/high/ctrlack_internal , 
        \I1/high/nlocalcd , \I1/high/U4/U28/U1/clr , \I1/high/U4/U28/U1/set , 
        \I1/high/U1/Z , \I1/high/U1664/y[0] , \I1/high/U1664/y[1] , 
        \I1/high/U1664/x[1] , \I1/high/U1664/x[3] , \I1/high/U1664/x[2] , 
        \I1/high/U1664/x[0] , \I1/high/U1664/U28/Z , \I1/high/U1664/U32/Z , 
        \I1/high/U1664/U29/Z , \I1/high/U1664/U33/Z , \I1/high/U1664/U30/Z , 
        \I1/high/U1664/U31/Z , \I1/high/U1664/U37/Z , \I1/high/U1669/nr , 
        \I1/high/U1669/nd , \I1/high/U1669/n2 , n1, n2, n3, n4, n5, n6, n7, n8;
    nand2_1 \U3/U5  ( .x(pullreq), .a(net30), .b(net31) );
    nor2_1 \I0/U3/U5  ( .x(net30), .a(\I0/net32 ), .b(\I0/net33 ) );
    buf_2 \I0/low/U1653  ( .x(\I0/low/latch ), .a(\I0/net32 ) );
    nor2_1 \I0/low/U264/U5  ( .x(\I0/low/nlocalcd ), .a(reset), .b(
        \I0/low/localcd ) );
    nor2_1 \I0/low/U1659_0_/U5  ( .x(\I0/low/ncd[0] ), .a(ol[0]), .b(oh[0]) );
    nor2_1 \I0/low/U1659_1_/U5  ( .x(\I0/low/ncd[1] ), .a(ol[1]), .b(oh[1]) );
    nor2_1 \I0/low/U1659_2_/U5  ( .x(\I0/low/ncd[2] ), .a(ol[2]), .b(oh[2]) );
    nor2_1 \I0/low/U1659_3_/U5  ( .x(\I0/low/ncd[3] ), .a(ol[3]), .b(oh[3]) );
    nor2_1 \I0/low/U1659_4_/U5  ( .x(\I0/low/ncd[4] ), .a(ol[4]), .b(oh[4]) );
    nor2_1 \I0/low/U1659_5_/U5  ( .x(\I0/low/ncd[5] ), .a(ol[5]), .b(oh[5]) );
    nor2_1 \I0/low/U1659_6_/U5  ( .x(\I0/low/ncd[6] ), .a(ol[6]), .b(oh[6]) );
    nor2_1 \I0/low/U1659_7_/U5  ( .x(\I0/low/ncd[7] ), .a(ol[7]), .b(oh[7]) );
    nor2_1 \I0/low/U3/U5  ( .x(\I0/low/ctrlack_internal ), .a(\I0/low/acb ), 
        .b(\I0/low/ba ) );
    buf_2 \I0/low/U1665/U7  ( .x(\I0/low/driveh ), .a(\I0/net20 ) );
    buf_2 \I0/low/U1666/U7  ( .x(\I0/low/drivel ), .a(\I0/net20 ) );
    ao23_1 \I0/low/U1658_0_/U21/U1/U1  ( .x(ol[0]), .a(\I0/low/driveh ), .b(ol
        [0]), .c(n1), .d(pull_l[0]), .e(n2) );
    ao23_1 \I0/low/U1658_1_/U21/U1/U1  ( .x(ol[1]), .a(\I0/low/drivel ), .b(ol
        [1]), .c(\I0/low/driveh ), .d(pull_l[1]), .e(n2) );
    ao23_1 \I0/low/U1658_2_/U21/U1/U1  ( .x(ol[2]), .a(\I0/low/drivel ), .b(ol
        [2]), .c(\I0/low/driveh ), .d(pull_l[2]), .e(n2) );
    ao23_1 \I0/low/U1658_3_/U21/U1/U1  ( .x(ol[3]), .a(\I0/low/driveh ), .b(ol
        [3]), .c(\I0/low/drivel ), .d(pull_l[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_4_/U21/U1/U1  ( .x(ol[4]), .a(n1), .b(ol[4]), .c(
        \I0/low/drivel ), .d(pull_l[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_5_/U21/U1/U1  ( .x(ol[5]), .a(\I0/low/driveh ), .b(ol
        [5]), .c(n1), .d(pull_l[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_6_/U21/U1/U1  ( .x(ol[6]), .a(\I0/low/drivel ), .b(ol
        [6]), .c(\I0/low/driveh ), .d(pull_l[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_7_/U21/U1/U1  ( .x(ol[7]), .a(n1), .b(ol[7]), .c(n1), 
        .d(pull_l[7]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_0_/U21/U1/U1  ( .x(oh[0]), .a(\I0/low/driveh ), .b(oh
        [0]), .c(n1), .d(pull_h[0]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_1_/U21/U1/U1  ( .x(oh[1]), .a(n1), .b(oh[1]), .c(
        \I0/low/drivel ), .d(pull_h[1]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_2_/U21/U1/U1  ( .x(oh[2]), .a(\I0/low/drivel ), .b(oh
        [2]), .c(\I0/low/drivel ), .d(pull_h[2]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_3_/U21/U1/U1  ( .x(oh[3]), .a(n1), .b(oh[3]), .c(
        \I0/low/driveh ), .d(pull_h[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_4_/U21/U1/U1  ( .x(oh[4]), .a(n1), .b(oh[4]), .c(n1), 
        .d(pull_h[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_5_/U21/U1/U1  ( .x(oh[5]), .a(\I0/low/drivel ), .b(oh
        [5]), .c(n1), .d(pull_h[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_6_/U21/U1/U1  ( .x(oh[6]), .a(\I0/low/drivel ), .b(oh
        [6]), .c(\I0/low/driveh ), .d(pull_h[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_7_/U21/U1/U1  ( .x(oh[7]), .a(\I0/low/driveh ), .b(oh
        [7]), .c(\I0/low/drivel ), .d(pull_h[7]), .e(\I0/low/latch ) );
    aoai211_1 \I0/low/U4/U28/U1/U1  ( .x(\I0/low/U4/U28/U1/clr ), .a(
        \I0/net20 ), .b(\I0/low/acb ), .c(\I0/low/nlocalcd ), .d(\I0/net32 )
         );
    nand3_1 \I0/low/U4/U28/U1/U2  ( .x(\I0/low/U4/U28/U1/set ), .a(
        \I0/low/nlocalcd ), .b(\I0/net20 ), .c(\I0/low/acb ) );
    nand2_2 \I0/low/U4/U28/U1/U3  ( .x(\I0/net32 ), .a(\I0/low/U4/U28/U1/clr ), 
        .b(\I0/low/U4/U28/U1/set ) );
    oai21_1 \I0/low/U1/U30/U1/U1  ( .x(\I0/low/acb ), .a(\I0/low/U1/Z ), .b(
        \I0/low/ba ), .c(\I0/net20 ) );
    inv_1 \I0/low/U1/U30/U1/U2  ( .x(\I0/low/U1/Z ), .a(\I0/low/acb ) );
    ao222_1 \I0/low/U5/U18/U1/U1  ( .x(\I0/low/ba ), .a(\I0/low/latch ), .b(
        pullcd), .c(\I0/low/latch ), .d(\I0/low/ba ), .e(pullcd), .f(
        \I0/low/ba ) );
    aoi222_1 \I0/low/U1664/U28/U30/U1  ( .x(\I0/low/U1664/x[3] ), .a(
        \I0/low/ncd[7] ), .b(\I0/low/ncd[6] ), .c(\I0/low/ncd[7] ), .d(
        \I0/low/U1664/U28/Z ), .e(\I0/low/ncd[6] ), .f(\I0/low/U1664/U28/Z )
         );
    inv_1 \I0/low/U1664/U28/U30/Uinv  ( .x(\I0/low/U1664/U28/Z ), .a(
        \I0/low/U1664/x[3] ) );
    aoi222_1 \I0/low/U1664/U32/U30/U1  ( .x(\I0/low/U1664/x[0] ), .a(
        \I0/low/ncd[1] ), .b(\I0/low/ncd[0] ), .c(\I0/low/ncd[1] ), .d(
        \I0/low/U1664/U32/Z ), .e(\I0/low/ncd[0] ), .f(\I0/low/U1664/U32/Z )
         );
    inv_1 \I0/low/U1664/U32/U30/Uinv  ( .x(\I0/low/U1664/U32/Z ), .a(
        \I0/low/U1664/x[0] ) );
    aoi222_1 \I0/low/U1664/U29/U30/U1  ( .x(\I0/low/U1664/x[2] ), .a(
        \I0/low/ncd[5] ), .b(\I0/low/ncd[4] ), .c(\I0/low/ncd[5] ), .d(
        \I0/low/U1664/U29/Z ), .e(\I0/low/ncd[4] ), .f(\I0/low/U1664/U29/Z )
         );
    inv_1 \I0/low/U1664/U29/U30/Uinv  ( .x(\I0/low/U1664/U29/Z ), .a(
        \I0/low/U1664/x[2] ) );
    aoi222_1 \I0/low/U1664/U33/U30/U1  ( .x(\I0/low/U1664/y[0] ), .a(
        \I0/low/U1664/x[1] ), .b(\I0/low/U1664/x[0] ), .c(\I0/low/U1664/x[1] ), 
        .d(\I0/low/U1664/U33/Z ), .e(\I0/low/U1664/x[0] ), .f(
        \I0/low/U1664/U33/Z ) );
    inv_1 \I0/low/U1664/U33/U30/Uinv  ( .x(\I0/low/U1664/U33/Z ), .a(
        \I0/low/U1664/y[0] ) );
    aoi222_1 \I0/low/U1664/U30/U30/U1  ( .x(\I0/low/U1664/y[1] ), .a(
        \I0/low/U1664/x[3] ), .b(\I0/low/U1664/x[2] ), .c(\I0/low/U1664/x[3] ), 
        .d(\I0/low/U1664/U30/Z ), .e(\I0/low/U1664/x[2] ), .f(
        \I0/low/U1664/U30/Z ) );
    inv_1 \I0/low/U1664/U30/U30/Uinv  ( .x(\I0/low/U1664/U30/Z ), .a(
        \I0/low/U1664/y[1] ) );
    aoi222_1 \I0/low/U1664/U31/U30/U1  ( .x(\I0/low/U1664/x[1] ), .a(
        \I0/low/ncd[3] ), .b(\I0/low/ncd[2] ), .c(\I0/low/ncd[3] ), .d(
        \I0/low/U1664/U31/Z ), .e(\I0/low/ncd[2] ), .f(\I0/low/U1664/U31/Z )
         );
    inv_1 \I0/low/U1664/U31/U30/Uinv  ( .x(\I0/low/U1664/U31/Z ), .a(
        \I0/low/U1664/x[1] ) );
    aoi222_1 \I0/low/U1664/U37/U30/U1  ( .x(\I0/low/localcd ), .a(
        \I0/low/U1664/y[0] ), .b(\I0/low/U1664/y[1] ), .c(\I0/low/U1664/y[0] ), 
        .d(\I0/low/U1664/U37/Z ), .e(\I0/low/U1664/y[1] ), .f(
        \I0/low/U1664/U37/Z ) );
    inv_1 \I0/low/U1664/U37/U30/Uinv  ( .x(\I0/low/U1664/U37/Z ), .a(
        \I0/low/localcd ) );
    nor3_1 \I0/low/U1669/Unr  ( .x(\I0/low/U1669/nr ), .a(
        \I0/low/ctrlack_internal ), .b(n1), .c(\I0/low/driveh ) );
    nand3_1 \I0/low/U1669/Und  ( .x(\I0/low/U1669/nd ), .a(
        \I0/low/ctrlack_internal ), .b(\I0/low/drivel ), .c(\I0/low/driveh )
         );
    oa21_1 \I0/low/U1669/U1  ( .x(\I0/low/U1669/n2 ), .a(\I0/low/U1669/n2 ), 
        .b(\I0/low/U1669/nr ), .c(\I0/low/U1669/nd ) );
    inv_2 \I0/low/U1669/U3  ( .x(ctrlack), .a(\I0/low/U1669/n2 ) );
    buf_2 \I0/high/U1653  ( .x(\I0/high/latch ), .a(\I0/net33 ) );
    nor2_1 \I0/high/U264/U5  ( .x(\I0/high/nlocalcd ), .a(reset), .b(
        \I0/high/localcd ) );
    nor2_1 \I0/high/U1659_0_/U5  ( .x(\I0/high/ncd[0] ), .a(ol[8]), .b(oh[8])
         );
    nor2_1 \I0/high/U1659_1_/U5  ( .x(\I0/high/ncd[1] ), .a(ol[9]), .b(oh[9])
         );
    nor2_1 \I0/high/U1659_2_/U5  ( .x(\I0/high/ncd[2] ), .a(ol[10]), .b(oh[10]
        ) );
    nor2_1 \I0/high/U1659_3_/U5  ( .x(\I0/high/ncd[3] ), .a(ol[11]), .b(oh[11]
        ) );
    nor2_1 \I0/high/U1659_4_/U5  ( .x(\I0/high/ncd[4] ), .a(ol[12]), .b(oh[12]
        ) );
    nor2_1 \I0/high/U1659_5_/U5  ( .x(\I0/high/ncd[5] ), .a(ol[13]), .b(oh[13]
        ) );
    nor2_1 \I0/high/U1659_6_/U5  ( .x(\I0/high/ncd[6] ), .a(ol[14]), .b(oh[14]
        ) );
    nor2_1 \I0/high/U1659_7_/U5  ( .x(\I0/high/ncd[7] ), .a(ol[15]), .b(oh[15]
        ) );
    nor2_1 \I0/high/U3/U5  ( .x(\I0/high/ctrlack_internal ), .a(\I0/high/acb ), 
        .b(\I0/high/ba ) );
    buf_2 \I0/high/U1665/U7  ( .x(\I0/high/driveh ), .a(net17) );
    buf_2 \I0/high/U1666/U7  ( .x(\I0/high/drivel ), .a(net17) );
    ao23_1 \I0/high/U1658_0_/U21/U1/U1  ( .x(ol[8]), .a(\I0/high/driveh ), .b(
        ol[8]), .c(n3), .d(pull_l[0]), .e(n4) );
    ao23_1 \I0/high/U1658_1_/U21/U1/U1  ( .x(ol[9]), .a(\I0/high/drivel ), .b(
        ol[9]), .c(\I0/high/driveh ), .d(pull_l[1]), .e(n4) );
    ao23_1 \I0/high/U1658_2_/U21/U1/U1  ( .x(ol[10]), .a(\I0/high/drivel ), 
        .b(ol[10]), .c(\I0/high/driveh ), .d(pull_l[2]), .e(n4) );
    ao23_1 \I0/high/U1658_3_/U21/U1/U1  ( .x(ol[11]), .a(\I0/high/driveh ), 
        .b(ol[11]), .c(\I0/high/drivel ), .d(pull_l[3]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_4_/U21/U1/U1  ( .x(ol[12]), .a(n3), .b(ol[12]), .c(
        \I0/high/drivel ), .d(pull_l[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_5_/U21/U1/U1  ( .x(ol[13]), .a(\I0/high/driveh ), 
        .b(ol[13]), .c(n3), .d(pull_l[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_6_/U21/U1/U1  ( .x(ol[14]), .a(\I0/high/drivel ), 
        .b(ol[14]), .c(\I0/high/driveh ), .d(pull_l[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_7_/U21/U1/U1  ( .x(ol[15]), .a(n3), .b(ol[15]), .c(
        n3), .d(pull_l[7]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_0_/U21/U1/U1  ( .x(oh[8]), .a(\I0/high/driveh ), .b(
        oh[8]), .c(n3), .d(pull_h[0]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_1_/U21/U1/U1  ( .x(oh[9]), .a(n3), .b(oh[9]), .c(
        \I0/high/drivel ), .d(pull_h[1]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_2_/U21/U1/U1  ( .x(oh[10]), .a(\I0/high/drivel ), 
        .b(oh[10]), .c(\I0/high/drivel ), .d(pull_h[2]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_3_/U21/U1/U1  ( .x(oh[11]), .a(n3), .b(oh[11]), .c(
        \I0/high/driveh ), .d(pull_h[3]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_4_/U21/U1/U1  ( .x(oh[12]), .a(n3), .b(oh[12]), .c(
        n3), .d(pull_h[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_5_/U21/U1/U1  ( .x(oh[13]), .a(\I0/high/drivel ), 
        .b(oh[13]), .c(n3), .d(pull_h[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_6_/U21/U1/U1  ( .x(oh[14]), .a(\I0/high/drivel ), 
        .b(oh[14]), .c(\I0/high/driveh ), .d(pull_h[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_7_/U21/U1/U1  ( .x(oh[15]), .a(\I0/high/driveh ), 
        .b(oh[15]), .c(\I0/high/drivel ), .d(pull_h[7]), .e(\I0/high/latch )
         );
    aoai211_1 \I0/high/U4/U28/U1/U1  ( .x(\I0/high/U4/U28/U1/clr ), .a(net17), 
        .b(\I0/high/acb ), .c(\I0/high/nlocalcd ), .d(\I0/net33 ) );
    nand3_1 \I0/high/U4/U28/U1/U2  ( .x(\I0/high/U4/U28/U1/set ), .a(
        \I0/high/nlocalcd ), .b(net17), .c(\I0/high/acb ) );
    nand2_2 \I0/high/U4/U28/U1/U3  ( .x(\I0/net33 ), .a(
        \I0/high/U4/U28/U1/clr ), .b(\I0/high/U4/U28/U1/set ) );
    oai21_1 \I0/high/U1/U30/U1/U1  ( .x(\I0/high/acb ), .a(\I0/high/U1/Z ), 
        .b(\I0/high/ba ), .c(net17) );
    inv_1 \I0/high/U1/U30/U1/U2  ( .x(\I0/high/U1/Z ), .a(\I0/high/acb ) );
    ao222_1 \I0/high/U5/U18/U1/U1  ( .x(\I0/high/ba ), .a(\I0/high/latch ), 
        .b(pullcd), .c(\I0/high/latch ), .d(\I0/high/ba ), .e(pullcd), .f(
        \I0/high/ba ) );
    aoi222_1 \I0/high/U1664/U28/U30/U1  ( .x(\I0/high/U1664/x[3] ), .a(
        \I0/high/ncd[7] ), .b(\I0/high/ncd[6] ), .c(\I0/high/ncd[7] ), .d(
        \I0/high/U1664/U28/Z ), .e(\I0/high/ncd[6] ), .f(\I0/high/U1664/U28/Z 
        ) );
    inv_1 \I0/high/U1664/U28/U30/Uinv  ( .x(\I0/high/U1664/U28/Z ), .a(
        \I0/high/U1664/x[3] ) );
    aoi222_1 \I0/high/U1664/U32/U30/U1  ( .x(\I0/high/U1664/x[0] ), .a(
        \I0/high/ncd[1] ), .b(\I0/high/ncd[0] ), .c(\I0/high/ncd[1] ), .d(
        \I0/high/U1664/U32/Z ), .e(\I0/high/ncd[0] ), .f(\I0/high/U1664/U32/Z 
        ) );
    inv_1 \I0/high/U1664/U32/U30/Uinv  ( .x(\I0/high/U1664/U32/Z ), .a(
        \I0/high/U1664/x[0] ) );
    aoi222_1 \I0/high/U1664/U29/U30/U1  ( .x(\I0/high/U1664/x[2] ), .a(
        \I0/high/ncd[5] ), .b(\I0/high/ncd[4] ), .c(\I0/high/ncd[5] ), .d(
        \I0/high/U1664/U29/Z ), .e(\I0/high/ncd[4] ), .f(\I0/high/U1664/U29/Z 
        ) );
    inv_1 \I0/high/U1664/U29/U30/Uinv  ( .x(\I0/high/U1664/U29/Z ), .a(
        \I0/high/U1664/x[2] ) );
    aoi222_1 \I0/high/U1664/U33/U30/U1  ( .x(\I0/high/U1664/y[0] ), .a(
        \I0/high/U1664/x[1] ), .b(\I0/high/U1664/x[0] ), .c(
        \I0/high/U1664/x[1] ), .d(\I0/high/U1664/U33/Z ), .e(
        \I0/high/U1664/x[0] ), .f(\I0/high/U1664/U33/Z ) );
    inv_1 \I0/high/U1664/U33/U30/Uinv  ( .x(\I0/high/U1664/U33/Z ), .a(
        \I0/high/U1664/y[0] ) );
    aoi222_1 \I0/high/U1664/U30/U30/U1  ( .x(\I0/high/U1664/y[1] ), .a(
        \I0/high/U1664/x[3] ), .b(\I0/high/U1664/x[2] ), .c(
        \I0/high/U1664/x[3] ), .d(\I0/high/U1664/U30/Z ), .e(
        \I0/high/U1664/x[2] ), .f(\I0/high/U1664/U30/Z ) );
    inv_1 \I0/high/U1664/U30/U30/Uinv  ( .x(\I0/high/U1664/U30/Z ), .a(
        \I0/high/U1664/y[1] ) );
    aoi222_1 \I0/high/U1664/U31/U30/U1  ( .x(\I0/high/U1664/x[1] ), .a(
        \I0/high/ncd[3] ), .b(\I0/high/ncd[2] ), .c(\I0/high/ncd[3] ), .d(
        \I0/high/U1664/U31/Z ), .e(\I0/high/ncd[2] ), .f(\I0/high/U1664/U31/Z 
        ) );
    inv_1 \I0/high/U1664/U31/U30/Uinv  ( .x(\I0/high/U1664/U31/Z ), .a(
        \I0/high/U1664/x[1] ) );
    aoi222_1 \I0/high/U1664/U37/U30/U1  ( .x(\I0/high/localcd ), .a(
        \I0/high/U1664/y[0] ), .b(\I0/high/U1664/y[1] ), .c(
        \I0/high/U1664/y[0] ), .d(\I0/high/U1664/U37/Z ), .e(
        \I0/high/U1664/y[1] ), .f(\I0/high/U1664/U37/Z ) );
    inv_1 \I0/high/U1664/U37/U30/Uinv  ( .x(\I0/high/U1664/U37/Z ), .a(
        \I0/high/localcd ) );
    nor3_1 \I0/high/U1669/Unr  ( .x(\I0/high/U1669/nr ), .a(
        \I0/high/ctrlack_internal ), .b(n3), .c(\I0/high/driveh ) );
    nand3_1 \I0/high/U1669/Und  ( .x(\I0/high/U1669/nd ), .a(
        \I0/high/ctrlack_internal ), .b(\I0/high/drivel ), .c(\I0/high/driveh 
        ) );
    oa21_1 \I0/high/U1669/U1  ( .x(\I0/high/U1669/n2 ), .a(\I0/high/U1669/n2 ), 
        .b(\I0/high/U1669/nr ), .c(\I0/high/U1669/nd ) );
    inv_2 \I0/high/U1669/U3  ( .x(\I0/net20 ), .a(\I0/high/U1669/n2 ) );
    nor2_1 \I1/U3/U5  ( .x(net31), .a(\I1/net32 ), .b(\I1/net33 ) );
    buf_2 \I1/low/U1653  ( .x(\I1/low/latch ), .a(\I1/net32 ) );
    nor2_1 \I1/low/U264/U5  ( .x(\I1/low/nlocalcd ), .a(reset), .b(
        \I1/low/localcd ) );
    nor2_1 \I1/low/U1659_0_/U5  ( .x(\I1/low/ncd[0] ), .a(ol[16]), .b(oh[16])
         );
    nor2_1 \I1/low/U1659_1_/U5  ( .x(\I1/low/ncd[1] ), .a(ol[17]), .b(oh[17])
         );
    nor2_1 \I1/low/U1659_2_/U5  ( .x(\I1/low/ncd[2] ), .a(ol[18]), .b(oh[18])
         );
    nor2_1 \I1/low/U1659_3_/U5  ( .x(\I1/low/ncd[3] ), .a(ol[19]), .b(oh[19])
         );
    nor2_1 \I1/low/U1659_4_/U5  ( .x(\I1/low/ncd[4] ), .a(ol[20]), .b(oh[20])
         );
    nor2_1 \I1/low/U1659_5_/U5  ( .x(\I1/low/ncd[5] ), .a(ol[21]), .b(oh[21])
         );
    nor2_1 \I1/low/U1659_6_/U5  ( .x(\I1/low/ncd[6] ), .a(ol[22]), .b(oh[22])
         );
    nor2_1 \I1/low/U1659_7_/U5  ( .x(\I1/low/ncd[7] ), .a(ol[23]), .b(oh[23])
         );
    nor2_1 \I1/low/U3/U5  ( .x(\I1/low/ctrlack_internal ), .a(\I1/low/acb ), 
        .b(\I1/low/ba ) );
    buf_2 \I1/low/U1665/U7  ( .x(\I1/low/driveh ), .a(\I1/net20 ) );
    buf_2 \I1/low/U1666/U7  ( .x(\I1/low/drivel ), .a(\I1/net20 ) );
    ao23_1 \I1/low/U1658_0_/U21/U1/U1  ( .x(ol[16]), .a(\I1/low/driveh ), .b(
        ol[16]), .c(n5), .d(pull_l[0]), .e(n6) );
    ao23_1 \I1/low/U1658_1_/U21/U1/U1  ( .x(ol[17]), .a(\I1/low/drivel ), .b(
        ol[17]), .c(\I1/low/driveh ), .d(pull_l[1]), .e(n6) );
    ao23_1 \I1/low/U1658_2_/U21/U1/U1  ( .x(ol[18]), .a(\I1/low/drivel ), .b(
        ol[18]), .c(\I1/low/driveh ), .d(pull_l[2]), .e(n6) );
    ao23_1 \I1/low/U1658_3_/U21/U1/U1  ( .x(ol[19]), .a(\I1/low/driveh ), .b(
        ol[19]), .c(\I1/low/drivel ), .d(pull_l[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_4_/U21/U1/U1  ( .x(ol[20]), .a(n5), .b(ol[20]), .c(
        \I1/low/drivel ), .d(pull_l[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_5_/U21/U1/U1  ( .x(ol[21]), .a(\I1/low/driveh ), .b(
        ol[21]), .c(n5), .d(pull_l[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_6_/U21/U1/U1  ( .x(ol[22]), .a(\I1/low/drivel ), .b(
        ol[22]), .c(\I1/low/driveh ), .d(pull_l[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_7_/U21/U1/U1  ( .x(ol[23]), .a(n5), .b(ol[23]), .c(n5
        ), .d(pull_l[7]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_0_/U21/U1/U1  ( .x(oh[16]), .a(\I1/low/driveh ), .b(
        oh[16]), .c(n5), .d(pull_h[0]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_1_/U21/U1/U1  ( .x(oh[17]), .a(n5), .b(oh[17]), .c(
        \I1/low/drivel ), .d(pull_h[1]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_2_/U21/U1/U1  ( .x(oh[18]), .a(\I1/low/drivel ), .b(
        oh[18]), .c(\I1/low/drivel ), .d(pull_h[2]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_3_/U21/U1/U1  ( .x(oh[19]), .a(n5), .b(oh[19]), .c(
        \I1/low/driveh ), .d(pull_h[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_4_/U21/U1/U1  ( .x(oh[20]), .a(n5), .b(oh[20]), .c(n5
        ), .d(pull_h[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_5_/U21/U1/U1  ( .x(oh[21]), .a(\I1/low/drivel ), .b(
        oh[21]), .c(n5), .d(pull_h[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_6_/U21/U1/U1  ( .x(oh[22]), .a(\I1/low/drivel ), .b(
        oh[22]), .c(\I1/low/driveh ), .d(pull_h[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_7_/U21/U1/U1  ( .x(oh[23]), .a(\I1/low/driveh ), .b(
        oh[23]), .c(\I1/low/drivel ), .d(pull_h[7]), .e(\I1/low/latch ) );
    aoai211_1 \I1/low/U4/U28/U1/U1  ( .x(\I1/low/U4/U28/U1/clr ), .a(
        \I1/net20 ), .b(\I1/low/acb ), .c(\I1/low/nlocalcd ), .d(\I1/net32 )
         );
    nand3_1 \I1/low/U4/U28/U1/U2  ( .x(\I1/low/U4/U28/U1/set ), .a(
        \I1/low/nlocalcd ), .b(\I1/net20 ), .c(\I1/low/acb ) );
    nand2_2 \I1/low/U4/U28/U1/U3  ( .x(\I1/net32 ), .a(\I1/low/U4/U28/U1/clr ), 
        .b(\I1/low/U4/U28/U1/set ) );
    oai21_1 \I1/low/U1/U30/U1/U1  ( .x(\I1/low/acb ), .a(\I1/low/U1/Z ), .b(
        \I1/low/ba ), .c(\I1/net20 ) );
    inv_1 \I1/low/U1/U30/U1/U2  ( .x(\I1/low/U1/Z ), .a(\I1/low/acb ) );
    ao222_1 \I1/low/U5/U18/U1/U1  ( .x(\I1/low/ba ), .a(\I1/low/latch ), .b(
        pullcd), .c(\I1/low/latch ), .d(\I1/low/ba ), .e(pullcd), .f(
        \I1/low/ba ) );
    aoi222_1 \I1/low/U1664/U28/U30/U1  ( .x(\I1/low/U1664/x[3] ), .a(
        \I1/low/ncd[7] ), .b(\I1/low/ncd[6] ), .c(\I1/low/ncd[7] ), .d(
        \I1/low/U1664/U28/Z ), .e(\I1/low/ncd[6] ), .f(\I1/low/U1664/U28/Z )
         );
    inv_1 \I1/low/U1664/U28/U30/Uinv  ( .x(\I1/low/U1664/U28/Z ), .a(
        \I1/low/U1664/x[3] ) );
    aoi222_1 \I1/low/U1664/U32/U30/U1  ( .x(\I1/low/U1664/x[0] ), .a(
        \I1/low/ncd[1] ), .b(\I1/low/ncd[0] ), .c(\I1/low/ncd[1] ), .d(
        \I1/low/U1664/U32/Z ), .e(\I1/low/ncd[0] ), .f(\I1/low/U1664/U32/Z )
         );
    inv_1 \I1/low/U1664/U32/U30/Uinv  ( .x(\I1/low/U1664/U32/Z ), .a(
        \I1/low/U1664/x[0] ) );
    aoi222_1 \I1/low/U1664/U29/U30/U1  ( .x(\I1/low/U1664/x[2] ), .a(
        \I1/low/ncd[5] ), .b(\I1/low/ncd[4] ), .c(\I1/low/ncd[5] ), .d(
        \I1/low/U1664/U29/Z ), .e(\I1/low/ncd[4] ), .f(\I1/low/U1664/U29/Z )
         );
    inv_1 \I1/low/U1664/U29/U30/Uinv  ( .x(\I1/low/U1664/U29/Z ), .a(
        \I1/low/U1664/x[2] ) );
    aoi222_1 \I1/low/U1664/U33/U30/U1  ( .x(\I1/low/U1664/y[0] ), .a(
        \I1/low/U1664/x[1] ), .b(\I1/low/U1664/x[0] ), .c(\I1/low/U1664/x[1] ), 
        .d(\I1/low/U1664/U33/Z ), .e(\I1/low/U1664/x[0] ), .f(
        \I1/low/U1664/U33/Z ) );
    inv_1 \I1/low/U1664/U33/U30/Uinv  ( .x(\I1/low/U1664/U33/Z ), .a(
        \I1/low/U1664/y[0] ) );
    aoi222_1 \I1/low/U1664/U30/U30/U1  ( .x(\I1/low/U1664/y[1] ), .a(
        \I1/low/U1664/x[3] ), .b(\I1/low/U1664/x[2] ), .c(\I1/low/U1664/x[3] ), 
        .d(\I1/low/U1664/U30/Z ), .e(\I1/low/U1664/x[2] ), .f(
        \I1/low/U1664/U30/Z ) );
    inv_1 \I1/low/U1664/U30/U30/Uinv  ( .x(\I1/low/U1664/U30/Z ), .a(
        \I1/low/U1664/y[1] ) );
    aoi222_1 \I1/low/U1664/U31/U30/U1  ( .x(\I1/low/U1664/x[1] ), .a(
        \I1/low/ncd[3] ), .b(\I1/low/ncd[2] ), .c(\I1/low/ncd[3] ), .d(
        \I1/low/U1664/U31/Z ), .e(\I1/low/ncd[2] ), .f(\I1/low/U1664/U31/Z )
         );
    inv_1 \I1/low/U1664/U31/U30/Uinv  ( .x(\I1/low/U1664/U31/Z ), .a(
        \I1/low/U1664/x[1] ) );
    aoi222_1 \I1/low/U1664/U37/U30/U1  ( .x(\I1/low/localcd ), .a(
        \I1/low/U1664/y[0] ), .b(\I1/low/U1664/y[1] ), .c(\I1/low/U1664/y[0] ), 
        .d(\I1/low/U1664/U37/Z ), .e(\I1/low/U1664/y[1] ), .f(
        \I1/low/U1664/U37/Z ) );
    inv_1 \I1/low/U1664/U37/U30/Uinv  ( .x(\I1/low/U1664/U37/Z ), .a(
        \I1/low/localcd ) );
    nor3_1 \I1/low/U1669/Unr  ( .x(\I1/low/U1669/nr ), .a(
        \I1/low/ctrlack_internal ), .b(n5), .c(\I1/low/driveh ) );
    nand3_1 \I1/low/U1669/Und  ( .x(\I1/low/U1669/nd ), .a(
        \I1/low/ctrlack_internal ), .b(\I1/low/drivel ), .c(\I1/low/driveh )
         );
    oa21_1 \I1/low/U1669/U1  ( .x(\I1/low/U1669/n2 ), .a(\I1/low/U1669/n2 ), 
        .b(\I1/low/U1669/nr ), .c(\I1/low/U1669/nd ) );
    inv_2 \I1/low/U1669/U3  ( .x(net17), .a(\I1/low/U1669/n2 ) );
    buf_2 \I1/high/U1653  ( .x(\I1/high/latch ), .a(\I1/net33 ) );
    nor2_1 \I1/high/U264/U5  ( .x(\I1/high/nlocalcd ), .a(reset), .b(
        \I1/high/localcd ) );
    nor2_1 \I1/high/U1659_0_/U5  ( .x(\I1/high/ncd[0] ), .a(ol[24]), .b(oh[24]
        ) );
    nor2_1 \I1/high/U1659_1_/U5  ( .x(\I1/high/ncd[1] ), .a(ol[25]), .b(oh[25]
        ) );
    nor2_1 \I1/high/U1659_2_/U5  ( .x(\I1/high/ncd[2] ), .a(ol[26]), .b(oh[26]
        ) );
    nor2_1 \I1/high/U1659_3_/U5  ( .x(\I1/high/ncd[3] ), .a(ol[27]), .b(oh[27]
        ) );
    nor2_1 \I1/high/U1659_4_/U5  ( .x(\I1/high/ncd[4] ), .a(ol[28]), .b(oh[28]
        ) );
    nor2_1 \I1/high/U1659_5_/U5  ( .x(\I1/high/ncd[5] ), .a(ol[29]), .b(oh[29]
        ) );
    nor2_1 \I1/high/U1659_6_/U5  ( .x(\I1/high/ncd[6] ), .a(ol[30]), .b(oh[30]
        ) );
    nor2_1 \I1/high/U1659_7_/U5  ( .x(\I1/high/ncd[7] ), .a(ol[31]), .b(oh[31]
        ) );
    nor2_1 \I1/high/U3/U5  ( .x(\I1/high/ctrlack_internal ), .a(\I1/high/acb ), 
        .b(\I1/high/ba ) );
    buf_2 \I1/high/U1665/U7  ( .x(\I1/high/driveh ), .a(ctrlreq) );
    buf_2 \I1/high/U1666/U7  ( .x(\I1/high/drivel ), .a(ctrlreq) );
    ao23_1 \I1/high/U1658_0_/U21/U1/U1  ( .x(ol[24]), .a(\I1/high/driveh ), 
        .b(ol[24]), .c(n7), .d(pull_l[0]), .e(n8) );
    ao23_1 \I1/high/U1658_1_/U21/U1/U1  ( .x(ol[25]), .a(\I1/high/drivel ), 
        .b(ol[25]), .c(\I1/high/driveh ), .d(pull_l[1]), .e(n8) );
    ao23_1 \I1/high/U1658_2_/U21/U1/U1  ( .x(ol[26]), .a(\I1/high/drivel ), 
        .b(ol[26]), .c(\I1/high/driveh ), .d(pull_l[2]), .e(n8) );
    ao23_1 \I1/high/U1658_3_/U21/U1/U1  ( .x(ol[27]), .a(\I1/high/driveh ), 
        .b(ol[27]), .c(\I1/high/drivel ), .d(pull_l[3]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1658_4_/U21/U1/U1  ( .x(ol[28]), .a(n7), .b(ol[28]), .c(
        \I1/high/drivel ), .d(pull_l[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_5_/U21/U1/U1  ( .x(ol[29]), .a(\I1/high/driveh ), 
        .b(ol[29]), .c(n7), .d(pull_l[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_6_/U21/U1/U1  ( .x(ol[30]), .a(\I1/high/drivel ), 
        .b(ol[30]), .c(\I1/high/driveh ), .d(pull_l[6]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1658_7_/U21/U1/U1  ( .x(ol[31]), .a(n7), .b(ol[31]), .c(
        n7), .d(pull_l[7]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_0_/U21/U1/U1  ( .x(oh[24]), .a(\I1/high/driveh ), 
        .b(oh[24]), .c(n7), .d(pull_h[0]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_1_/U21/U1/U1  ( .x(oh[25]), .a(n7), .b(oh[25]), .c(
        \I1/high/drivel ), .d(pull_h[1]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_2_/U21/U1/U1  ( .x(oh[26]), .a(\I1/high/drivel ), 
        .b(oh[26]), .c(\I1/high/drivel ), .d(pull_h[2]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1651_3_/U21/U1/U1  ( .x(oh[27]), .a(n7), .b(oh[27]), .c(
        \I1/high/driveh ), .d(pull_h[3]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_4_/U21/U1/U1  ( .x(oh[28]), .a(n7), .b(oh[28]), .c(
        n7), .d(pull_h[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_5_/U21/U1/U1  ( .x(oh[29]), .a(\I1/high/drivel ), 
        .b(oh[29]), .c(n7), .d(pull_h[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_6_/U21/U1/U1  ( .x(oh[30]), .a(\I1/high/drivel ), 
        .b(oh[30]), .c(\I1/high/driveh ), .d(pull_h[6]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1651_7_/U21/U1/U1  ( .x(oh[31]), .a(\I1/high/driveh ), 
        .b(oh[31]), .c(\I1/high/drivel ), .d(pull_h[7]), .e(\I1/high/latch )
         );
    aoai211_1 \I1/high/U4/U28/U1/U1  ( .x(\I1/high/U4/U28/U1/clr ), .a(ctrlreq
        ), .b(\I1/high/acb ), .c(\I1/high/nlocalcd ), .d(\I1/net33 ) );
    nand3_1 \I1/high/U4/U28/U1/U2  ( .x(\I1/high/U4/U28/U1/set ), .a(
        \I1/high/nlocalcd ), .b(ctrlreq), .c(\I1/high/acb ) );
    nand2_2 \I1/high/U4/U28/U1/U3  ( .x(\I1/net33 ), .a(
        \I1/high/U4/U28/U1/clr ), .b(\I1/high/U4/U28/U1/set ) );
    oai21_1 \I1/high/U1/U30/U1/U1  ( .x(\I1/high/acb ), .a(\I1/high/U1/Z ), 
        .b(\I1/high/ba ), .c(ctrlreq) );
    inv_1 \I1/high/U1/U30/U1/U2  ( .x(\I1/high/U1/Z ), .a(\I1/high/acb ) );
    ao222_1 \I1/high/U5/U18/U1/U1  ( .x(\I1/high/ba ), .a(\I1/high/latch ), 
        .b(pullcd), .c(\I1/high/latch ), .d(\I1/high/ba ), .e(pullcd), .f(
        \I1/high/ba ) );
    aoi222_1 \I1/high/U1664/U28/U30/U1  ( .x(\I1/high/U1664/x[3] ), .a(
        \I1/high/ncd[7] ), .b(\I1/high/ncd[6] ), .c(\I1/high/ncd[7] ), .d(
        \I1/high/U1664/U28/Z ), .e(\I1/high/ncd[6] ), .f(\I1/high/U1664/U28/Z 
        ) );
    inv_1 \I1/high/U1664/U28/U30/Uinv  ( .x(\I1/high/U1664/U28/Z ), .a(
        \I1/high/U1664/x[3] ) );
    aoi222_1 \I1/high/U1664/U32/U30/U1  ( .x(\I1/high/U1664/x[0] ), .a(
        \I1/high/ncd[1] ), .b(\I1/high/ncd[0] ), .c(\I1/high/ncd[1] ), .d(
        \I1/high/U1664/U32/Z ), .e(\I1/high/ncd[0] ), .f(\I1/high/U1664/U32/Z 
        ) );
    inv_1 \I1/high/U1664/U32/U30/Uinv  ( .x(\I1/high/U1664/U32/Z ), .a(
        \I1/high/U1664/x[0] ) );
    aoi222_1 \I1/high/U1664/U29/U30/U1  ( .x(\I1/high/U1664/x[2] ), .a(
        \I1/high/ncd[5] ), .b(\I1/high/ncd[4] ), .c(\I1/high/ncd[5] ), .d(
        \I1/high/U1664/U29/Z ), .e(\I1/high/ncd[4] ), .f(\I1/high/U1664/U29/Z 
        ) );
    inv_1 \I1/high/U1664/U29/U30/Uinv  ( .x(\I1/high/U1664/U29/Z ), .a(
        \I1/high/U1664/x[2] ) );
    aoi222_1 \I1/high/U1664/U33/U30/U1  ( .x(\I1/high/U1664/y[0] ), .a(
        \I1/high/U1664/x[1] ), .b(\I1/high/U1664/x[0] ), .c(
        \I1/high/U1664/x[1] ), .d(\I1/high/U1664/U33/Z ), .e(
        \I1/high/U1664/x[0] ), .f(\I1/high/U1664/U33/Z ) );
    inv_1 \I1/high/U1664/U33/U30/Uinv  ( .x(\I1/high/U1664/U33/Z ), .a(
        \I1/high/U1664/y[0] ) );
    aoi222_1 \I1/high/U1664/U30/U30/U1  ( .x(\I1/high/U1664/y[1] ), .a(
        \I1/high/U1664/x[3] ), .b(\I1/high/U1664/x[2] ), .c(
        \I1/high/U1664/x[3] ), .d(\I1/high/U1664/U30/Z ), .e(
        \I1/high/U1664/x[2] ), .f(\I1/high/U1664/U30/Z ) );
    inv_1 \I1/high/U1664/U30/U30/Uinv  ( .x(\I1/high/U1664/U30/Z ), .a(
        \I1/high/U1664/y[1] ) );
    aoi222_1 \I1/high/U1664/U31/U30/U1  ( .x(\I1/high/U1664/x[1] ), .a(
        \I1/high/ncd[3] ), .b(\I1/high/ncd[2] ), .c(\I1/high/ncd[3] ), .d(
        \I1/high/U1664/U31/Z ), .e(\I1/high/ncd[2] ), .f(\I1/high/U1664/U31/Z 
        ) );
    inv_1 \I1/high/U1664/U31/U30/Uinv  ( .x(\I1/high/U1664/U31/Z ), .a(
        \I1/high/U1664/x[1] ) );
    aoi222_1 \I1/high/U1664/U37/U30/U1  ( .x(\I1/high/localcd ), .a(
        \I1/high/U1664/y[0] ), .b(\I1/high/U1664/y[1] ), .c(
        \I1/high/U1664/y[0] ), .d(\I1/high/U1664/U37/Z ), .e(
        \I1/high/U1664/y[1] ), .f(\I1/high/U1664/U37/Z ) );
    inv_1 \I1/high/U1664/U37/U30/Uinv  ( .x(\I1/high/U1664/U37/Z ), .a(
        \I1/high/localcd ) );
    nor3_1 \I1/high/U1669/Unr  ( .x(\I1/high/U1669/nr ), .a(
        \I1/high/ctrlack_internal ), .b(n7), .c(\I1/high/driveh ) );
    nand3_1 \I1/high/U1669/Und  ( .x(\I1/high/U1669/nd ), .a(
        \I1/high/ctrlack_internal ), .b(\I1/high/drivel ), .c(\I1/high/driveh 
        ) );
    oa21_1 \I1/high/U1669/U1  ( .x(\I1/high/U1669/n2 ), .a(\I1/high/U1669/n2 ), 
        .b(\I1/high/U1669/nr ), .c(\I1/high/U1669/nd ) );
    inv_2 \I1/high/U1669/U3  ( .x(\I1/net20 ), .a(\I1/high/U1669/n2 ) );
    buf_2 U1 ( .x(n1), .a(\I0/net20 ) );
    buf_1 U2 ( .x(n2), .a(\I0/low/latch ) );
    buf_2 U3 ( .x(n3), .a(net17) );
    buf_1 U4 ( .x(n4), .a(\I0/high/latch ) );
    buf_2 U5 ( .x(n5), .a(\I1/net20 ) );
    buf_1 U6 ( .x(n6), .a(\I1/low/latch ) );
    buf_2 U7 ( .x(n7), .a(ctrlreq) );
    buf_1 U8 ( .x(n8), .a(\I1/high/latch ) );
endmodule


module chain_irdemux_32new_1 ( ctrlack, oh, ol, pullreq, pull_h, pull_l, 
    pullcd, reset, ctrlreq );
output [31:0] oh;
output [31:0] ol;
input  [7:0] pull_h;
input  [7:0] pull_l;
input  pullcd, reset, ctrlreq;
output ctrlack, pullreq;
    wire net30, net31, net17, \I0/net20 , \I0/net33 , \I0/net32 , 
        \I0/low/drivel , \I0/low/driveh , \I0/low/localcd , \I0/low/ncd[7] , 
        \I0/low/ncd[6] , \I0/low/ncd[5] , \I0/low/ncd[4] , \I0/low/ncd[3] , 
        \I0/low/ncd[2] , \I0/low/ncd[1] , \I0/low/ncd[0] , \I0/low/ba , 
        \I0/low/latch , \I0/low/acb , \I0/low/ctrlack_internal , 
        \I0/low/nlocalcd , \I0/low/U4/U28/U1/clr , \I0/low/U4/U28/U1/set , 
        \I0/low/U1/Z , \I0/low/U1664/y[0] , \I0/low/U1664/y[1] , 
        \I0/low/U1664/x[1] , \I0/low/U1664/x[3] , \I0/low/U1664/x[2] , 
        \I0/low/U1664/x[0] , \I0/low/U1664/U28/Z , \I0/low/U1664/U32/Z , 
        \I0/low/U1664/U29/Z , \I0/low/U1664/U33/Z , \I0/low/U1664/U30/Z , 
        \I0/low/U1664/U31/Z , \I0/low/U1664/U37/Z , \I0/low/U1669/nr , 
        \I0/low/U1669/nd , \I0/low/U1669/n2 , \I0/high/drivel , 
        \I0/high/driveh , \I0/high/localcd , \I0/high/ncd[7] , 
        \I0/high/ncd[6] , \I0/high/ncd[5] , \I0/high/ncd[4] , \I0/high/ncd[3] , 
        \I0/high/ncd[2] , \I0/high/ncd[1] , \I0/high/ncd[0] , \I0/high/ba , 
        \I0/high/latch , \I0/high/acb , \I0/high/ctrlack_internal , 
        \I0/high/nlocalcd , \I0/high/U4/U28/U1/clr , \I0/high/U4/U28/U1/set , 
        \I0/high/U1/Z , \I0/high/U1664/y[0] , \I0/high/U1664/y[1] , 
        \I0/high/U1664/x[1] , \I0/high/U1664/x[3] , \I0/high/U1664/x[2] , 
        \I0/high/U1664/x[0] , \I0/high/U1664/U28/Z , \I0/high/U1664/U32/Z , 
        \I0/high/U1664/U29/Z , \I0/high/U1664/U33/Z , \I0/high/U1664/U30/Z , 
        \I0/high/U1664/U31/Z , \I0/high/U1664/U37/Z , \I0/high/U1669/nr , 
        \I0/high/U1669/nd , \I0/high/U1669/n2 , \I1/net20 , \I1/net33 , 
        \I1/net32 , \I1/low/drivel , \I1/low/driveh , \I1/low/localcd , 
        \I1/low/ncd[7] , \I1/low/ncd[6] , \I1/low/ncd[5] , \I1/low/ncd[4] , 
        \I1/low/ncd[3] , \I1/low/ncd[2] , \I1/low/ncd[1] , \I1/low/ncd[0] , 
        \I1/low/ba , \I1/low/latch , \I1/low/acb , \I1/low/ctrlack_internal , 
        \I1/low/nlocalcd , \I1/low/U4/U28/U1/clr , \I1/low/U4/U28/U1/set , 
        \I1/low/U1/Z , \I1/low/U1664/y[0] , \I1/low/U1664/y[1] , 
        \I1/low/U1664/x[1] , \I1/low/U1664/x[3] , \I1/low/U1664/x[2] , 
        \I1/low/U1664/x[0] , \I1/low/U1664/U28/Z , \I1/low/U1664/U32/Z , 
        \I1/low/U1664/U29/Z , \I1/low/U1664/U33/Z , \I1/low/U1664/U30/Z , 
        \I1/low/U1664/U31/Z , \I1/low/U1664/U37/Z , \I1/low/U1669/nr , 
        \I1/low/U1669/nd , \I1/low/U1669/n2 , \I1/high/localcd , 
        \I1/high/ncd[7] , \I1/high/ncd[6] , \I1/high/ncd[5] , \I1/high/ncd[4] , 
        \I1/high/ncd[3] , \I1/high/ncd[2] , \I1/high/ncd[1] , \I1/high/ncd[0] , 
        \I1/high/ba , \I1/high/latch , \I1/high/acb , 
        \I1/high/ctrlack_internal , \I1/high/nlocalcd , 
        \I1/high/U4/U28/U1/clr , \I1/high/U4/U28/U1/set , \I1/high/U1/Z , 
        \I1/high/U1664/y[0] , \I1/high/U1664/y[1] , \I1/high/U1664/x[1] , 
        \I1/high/U1664/x[3] , \I1/high/U1664/x[2] , \I1/high/U1664/x[0] , 
        \I1/high/U1664/U28/Z , \I1/high/U1664/U32/Z , \I1/high/U1664/U29/Z , 
        \I1/high/U1664/U33/Z , \I1/high/U1664/U30/Z , \I1/high/U1664/U31/Z , 
        \I1/high/U1664/U37/Z , \I1/high/U1669/nr , \I1/high/U1669/nd , 
        \I1/high/U1669/n2 , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
    nand2_1 \U3/U5  ( .x(pullreq), .a(net30), .b(net31) );
    nor2_1 \I0/U3/U5  ( .x(net30), .a(\I0/net32 ), .b(\I0/net33 ) );
    buf_2 \I0/low/U1653  ( .x(\I0/low/latch ), .a(\I0/net32 ) );
    nor2_1 \I0/low/U264/U5  ( .x(\I0/low/nlocalcd ), .a(reset), .b(
        \I0/low/localcd ) );
    nor2_1 \I0/low/U1659_0_/U5  ( .x(\I0/low/ncd[0] ), .a(ol[0]), .b(oh[0]) );
    nor2_1 \I0/low/U1659_1_/U5  ( .x(\I0/low/ncd[1] ), .a(ol[1]), .b(oh[1]) );
    nor2_1 \I0/low/U1659_2_/U5  ( .x(\I0/low/ncd[2] ), .a(ol[2]), .b(oh[2]) );
    nor2_1 \I0/low/U1659_3_/U5  ( .x(\I0/low/ncd[3] ), .a(ol[3]), .b(oh[3]) );
    nor2_1 \I0/low/U1659_4_/U5  ( .x(\I0/low/ncd[4] ), .a(ol[4]), .b(oh[4]) );
    nor2_1 \I0/low/U1659_5_/U5  ( .x(\I0/low/ncd[5] ), .a(ol[5]), .b(oh[5]) );
    nor2_1 \I0/low/U1659_6_/U5  ( .x(\I0/low/ncd[6] ), .a(ol[6]), .b(oh[6]) );
    nor2_1 \I0/low/U1659_7_/U5  ( .x(\I0/low/ncd[7] ), .a(ol[7]), .b(oh[7]) );
    nor2_1 \I0/low/U3/U5  ( .x(\I0/low/ctrlack_internal ), .a(\I0/low/acb ), 
        .b(\I0/low/ba ) );
    buf_2 \I0/low/U1665/U7  ( .x(\I0/low/driveh ), .a(\I0/net20 ) );
    buf_2 \I0/low/U1666/U7  ( .x(\I0/low/drivel ), .a(\I0/net20 ) );
    ao23_1 \I0/low/U1658_0_/U21/U1/U1  ( .x(ol[0]), .a(n12), .b(ol[0]), .c(
        \I0/low/drivel ), .d(pull_l[0]), .e(n11) );
    ao23_1 \I0/low/U1658_1_/U21/U1/U1  ( .x(ol[1]), .a(n12), .b(ol[1]), .c(
        \I0/low/driveh ), .d(pull_l[1]), .e(n11) );
    ao23_1 \I0/low/U1658_2_/U21/U1/U1  ( .x(ol[2]), .a(\I0/low/driveh ), .b(ol
        [2]), .c(n12), .d(pull_l[2]), .e(n11) );
    ao23_1 \I0/low/U1658_3_/U21/U1/U1  ( .x(ol[3]), .a(n12), .b(ol[3]), .c(
        \I0/low/driveh ), .d(pull_l[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_4_/U21/U1/U1  ( .x(ol[4]), .a(\I0/low/drivel ), .b(ol
        [4]), .c(n12), .d(pull_l[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_5_/U21/U1/U1  ( .x(ol[5]), .a(\I0/low/drivel ), .b(ol
        [5]), .c(n12), .d(pull_l[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_6_/U21/U1/U1  ( .x(ol[6]), .a(\I0/low/driveh ), .b(ol
        [6]), .c(\I0/low/drivel ), .d(pull_l[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_7_/U21/U1/U1  ( .x(ol[7]), .a(\I0/low/driveh ), .b(ol
        [7]), .c(\I0/low/driveh ), .d(pull_l[7]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_0_/U21/U1/U1  ( .x(oh[0]), .a(\I0/low/drivel ), .b(oh
        [0]), .c(n12), .d(pull_h[0]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_1_/U21/U1/U1  ( .x(oh[1]), .a(\I0/low/driveh ), .b(oh
        [1]), .c(\I0/low/drivel ), .d(pull_h[1]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_2_/U21/U1/U1  ( .x(oh[2]), .a(\I0/low/drivel ), .b(oh
        [2]), .c(\I0/low/drivel ), .d(pull_h[2]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_3_/U21/U1/U1  ( .x(oh[3]), .a(\I0/low/driveh ), .b(oh
        [3]), .c(\I0/low/driveh ), .d(pull_h[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_4_/U21/U1/U1  ( .x(oh[4]), .a(\I0/low/drivel ), .b(oh
        [4]), .c(\I0/low/driveh ), .d(pull_h[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_5_/U21/U1/U1  ( .x(oh[5]), .a(\I0/low/driveh ), .b(oh
        [5]), .c(n12), .d(pull_h[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_6_/U21/U1/U1  ( .x(oh[6]), .a(n12), .b(oh[6]), .c(
        \I0/low/drivel ), .d(pull_h[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_7_/U21/U1/U1  ( .x(oh[7]), .a(n12), .b(oh[7]), .c(n12
        ), .d(pull_h[7]), .e(\I0/low/latch ) );
    aoai211_1 \I0/low/U4/U28/U1/U1  ( .x(\I0/low/U4/U28/U1/clr ), .a(
        \I0/net20 ), .b(\I0/low/acb ), .c(\I0/low/nlocalcd ), .d(\I0/net32 )
         );
    nand3_1 \I0/low/U4/U28/U1/U2  ( .x(\I0/low/U4/U28/U1/set ), .a(
        \I0/low/nlocalcd ), .b(\I0/net20 ), .c(\I0/low/acb ) );
    nand2_2 \I0/low/U4/U28/U1/U3  ( .x(\I0/net32 ), .a(\I0/low/U4/U28/U1/clr ), 
        .b(\I0/low/U4/U28/U1/set ) );
    oai21_1 \I0/low/U1/U30/U1/U1  ( .x(\I0/low/acb ), .a(\I0/low/U1/Z ), .b(
        \I0/low/ba ), .c(\I0/net20 ) );
    inv_1 \I0/low/U1/U30/U1/U2  ( .x(\I0/low/U1/Z ), .a(\I0/low/acb ) );
    ao222_1 \I0/low/U5/U18/U1/U1  ( .x(\I0/low/ba ), .a(\I0/low/latch ), .b(
        pullcd), .c(\I0/low/latch ), .d(\I0/low/ba ), .e(pullcd), .f(
        \I0/low/ba ) );
    aoi222_1 \I0/low/U1664/U28/U30/U1  ( .x(\I0/low/U1664/x[3] ), .a(
        \I0/low/ncd[7] ), .b(\I0/low/ncd[6] ), .c(\I0/low/ncd[7] ), .d(
        \I0/low/U1664/U28/Z ), .e(\I0/low/ncd[6] ), .f(\I0/low/U1664/U28/Z )
         );
    inv_1 \I0/low/U1664/U28/U30/Uinv  ( .x(\I0/low/U1664/U28/Z ), .a(
        \I0/low/U1664/x[3] ) );
    aoi222_1 \I0/low/U1664/U32/U30/U1  ( .x(\I0/low/U1664/x[0] ), .a(
        \I0/low/ncd[1] ), .b(\I0/low/ncd[0] ), .c(\I0/low/ncd[1] ), .d(
        \I0/low/U1664/U32/Z ), .e(\I0/low/ncd[0] ), .f(\I0/low/U1664/U32/Z )
         );
    inv_1 \I0/low/U1664/U32/U30/Uinv  ( .x(\I0/low/U1664/U32/Z ), .a(
        \I0/low/U1664/x[0] ) );
    aoi222_1 \I0/low/U1664/U29/U30/U1  ( .x(\I0/low/U1664/x[2] ), .a(
        \I0/low/ncd[5] ), .b(\I0/low/ncd[4] ), .c(\I0/low/ncd[5] ), .d(
        \I0/low/U1664/U29/Z ), .e(\I0/low/ncd[4] ), .f(\I0/low/U1664/U29/Z )
         );
    inv_1 \I0/low/U1664/U29/U30/Uinv  ( .x(\I0/low/U1664/U29/Z ), .a(
        \I0/low/U1664/x[2] ) );
    aoi222_1 \I0/low/U1664/U33/U30/U1  ( .x(\I0/low/U1664/y[0] ), .a(
        \I0/low/U1664/x[1] ), .b(\I0/low/U1664/x[0] ), .c(\I0/low/U1664/x[1] ), 
        .d(\I0/low/U1664/U33/Z ), .e(\I0/low/U1664/x[0] ), .f(
        \I0/low/U1664/U33/Z ) );
    inv_1 \I0/low/U1664/U33/U30/Uinv  ( .x(\I0/low/U1664/U33/Z ), .a(
        \I0/low/U1664/y[0] ) );
    aoi222_1 \I0/low/U1664/U30/U30/U1  ( .x(\I0/low/U1664/y[1] ), .a(
        \I0/low/U1664/x[3] ), .b(\I0/low/U1664/x[2] ), .c(\I0/low/U1664/x[3] ), 
        .d(\I0/low/U1664/U30/Z ), .e(\I0/low/U1664/x[2] ), .f(
        \I0/low/U1664/U30/Z ) );
    inv_1 \I0/low/U1664/U30/U30/Uinv  ( .x(\I0/low/U1664/U30/Z ), .a(
        \I0/low/U1664/y[1] ) );
    aoi222_1 \I0/low/U1664/U31/U30/U1  ( .x(\I0/low/U1664/x[1] ), .a(
        \I0/low/ncd[3] ), .b(\I0/low/ncd[2] ), .c(\I0/low/ncd[3] ), .d(
        \I0/low/U1664/U31/Z ), .e(\I0/low/ncd[2] ), .f(\I0/low/U1664/U31/Z )
         );
    inv_1 \I0/low/U1664/U31/U30/Uinv  ( .x(\I0/low/U1664/U31/Z ), .a(
        \I0/low/U1664/x[1] ) );
    aoi222_1 \I0/low/U1664/U37/U30/U1  ( .x(\I0/low/localcd ), .a(
        \I0/low/U1664/y[0] ), .b(\I0/low/U1664/y[1] ), .c(\I0/low/U1664/y[0] ), 
        .d(\I0/low/U1664/U37/Z ), .e(\I0/low/U1664/y[1] ), .f(
        \I0/low/U1664/U37/Z ) );
    inv_1 \I0/low/U1664/U37/U30/Uinv  ( .x(\I0/low/U1664/U37/Z ), .a(
        \I0/low/localcd ) );
    nor3_1 \I0/low/U1669/Unr  ( .x(\I0/low/U1669/nr ), .a(
        \I0/low/ctrlack_internal ), .b(n12), .c(\I0/low/drivel ) );
    nand3_1 \I0/low/U1669/Und  ( .x(\I0/low/U1669/nd ), .a(
        \I0/low/ctrlack_internal ), .b(\I0/low/driveh ), .c(\I0/low/drivel )
         );
    oa21_1 \I0/low/U1669/U1  ( .x(\I0/low/U1669/n2 ), .a(\I0/low/U1669/n2 ), 
        .b(\I0/low/U1669/nr ), .c(\I0/low/U1669/nd ) );
    inv_2 \I0/low/U1669/U3  ( .x(ctrlack), .a(\I0/low/U1669/n2 ) );
    buf_2 \I0/high/U1653  ( .x(\I0/high/latch ), .a(\I0/net33 ) );
    nor2_1 \I0/high/U264/U5  ( .x(\I0/high/nlocalcd ), .a(reset), .b(
        \I0/high/localcd ) );
    nor2_1 \I0/high/U1659_0_/U5  ( .x(\I0/high/ncd[0] ), .a(ol[8]), .b(oh[8])
         );
    nor2_1 \I0/high/U1659_1_/U5  ( .x(\I0/high/ncd[1] ), .a(ol[9]), .b(oh[9])
         );
    nor2_1 \I0/high/U1659_2_/U5  ( .x(\I0/high/ncd[2] ), .a(ol[10]), .b(oh[10]
        ) );
    nor2_1 \I0/high/U1659_3_/U5  ( .x(\I0/high/ncd[3] ), .a(ol[11]), .b(oh[11]
        ) );
    nor2_1 \I0/high/U1659_4_/U5  ( .x(\I0/high/ncd[4] ), .a(ol[12]), .b(oh[12]
        ) );
    nor2_1 \I0/high/U1659_5_/U5  ( .x(\I0/high/ncd[5] ), .a(ol[13]), .b(oh[13]
        ) );
    nor2_1 \I0/high/U1659_6_/U5  ( .x(\I0/high/ncd[6] ), .a(ol[14]), .b(oh[14]
        ) );
    nor2_1 \I0/high/U1659_7_/U5  ( .x(\I0/high/ncd[7] ), .a(ol[15]), .b(oh[15]
        ) );
    nor2_1 \I0/high/U3/U5  ( .x(\I0/high/ctrlack_internal ), .a(\I0/high/acb ), 
        .b(\I0/high/ba ) );
    buf_2 \I0/high/U1665/U7  ( .x(\I0/high/driveh ), .a(net17) );
    buf_2 \I0/high/U1666/U7  ( .x(\I0/high/drivel ), .a(net17) );
    ao23_1 \I0/high/U1658_0_/U21/U1/U1  ( .x(ol[8]), .a(n10), .b(ol[8]), .c(
        \I0/high/drivel ), .d(pull_l[0]), .e(n9) );
    ao23_1 \I0/high/U1658_1_/U21/U1/U1  ( .x(ol[9]), .a(n10), .b(ol[9]), .c(
        \I0/high/driveh ), .d(pull_l[1]), .e(n9) );
    ao23_1 \I0/high/U1658_2_/U21/U1/U1  ( .x(ol[10]), .a(\I0/high/driveh ), 
        .b(ol[10]), .c(n10), .d(pull_l[2]), .e(n9) );
    ao23_1 \I0/high/U1658_3_/U21/U1/U1  ( .x(ol[11]), .a(n10), .b(ol[11]), .c(
        \I0/high/driveh ), .d(pull_l[3]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_4_/U21/U1/U1  ( .x(ol[12]), .a(\I0/high/drivel ), 
        .b(ol[12]), .c(n10), .d(pull_l[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_5_/U21/U1/U1  ( .x(ol[13]), .a(\I0/high/drivel ), 
        .b(ol[13]), .c(n10), .d(pull_l[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_6_/U21/U1/U1  ( .x(ol[14]), .a(\I0/high/driveh ), 
        .b(ol[14]), .c(\I0/high/drivel ), .d(pull_l[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_7_/U21/U1/U1  ( .x(ol[15]), .a(\I0/high/driveh ), 
        .b(ol[15]), .c(\I0/high/driveh ), .d(pull_l[7]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_0_/U21/U1/U1  ( .x(oh[8]), .a(\I0/high/drivel ), .b(
        oh[8]), .c(n10), .d(pull_h[0]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_1_/U21/U1/U1  ( .x(oh[9]), .a(\I0/high/driveh ), .b(
        oh[9]), .c(\I0/high/drivel ), .d(pull_h[1]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_2_/U21/U1/U1  ( .x(oh[10]), .a(\I0/high/drivel ), 
        .b(oh[10]), .c(\I0/high/drivel ), .d(pull_h[2]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_3_/U21/U1/U1  ( .x(oh[11]), .a(\I0/high/driveh ), 
        .b(oh[11]), .c(\I0/high/driveh ), .d(pull_h[3]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_4_/U21/U1/U1  ( .x(oh[12]), .a(\I0/high/drivel ), 
        .b(oh[12]), .c(\I0/high/driveh ), .d(pull_h[4]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_5_/U21/U1/U1  ( .x(oh[13]), .a(\I0/high/driveh ), 
        .b(oh[13]), .c(n10), .d(pull_h[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_6_/U21/U1/U1  ( .x(oh[14]), .a(n10), .b(oh[14]), .c(
        \I0/high/drivel ), .d(pull_h[6]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_7_/U21/U1/U1  ( .x(oh[15]), .a(n10), .b(oh[15]), .c(
        n10), .d(pull_h[7]), .e(\I0/high/latch ) );
    aoai211_1 \I0/high/U4/U28/U1/U1  ( .x(\I0/high/U4/U28/U1/clr ), .a(net17), 
        .b(\I0/high/acb ), .c(\I0/high/nlocalcd ), .d(\I0/net33 ) );
    nand3_1 \I0/high/U4/U28/U1/U2  ( .x(\I0/high/U4/U28/U1/set ), .a(
        \I0/high/nlocalcd ), .b(net17), .c(\I0/high/acb ) );
    nand2_2 \I0/high/U4/U28/U1/U3  ( .x(\I0/net33 ), .a(
        \I0/high/U4/U28/U1/clr ), .b(\I0/high/U4/U28/U1/set ) );
    oai21_1 \I0/high/U1/U30/U1/U1  ( .x(\I0/high/acb ), .a(\I0/high/U1/Z ), 
        .b(\I0/high/ba ), .c(net17) );
    inv_1 \I0/high/U1/U30/U1/U2  ( .x(\I0/high/U1/Z ), .a(\I0/high/acb ) );
    ao222_1 \I0/high/U5/U18/U1/U1  ( .x(\I0/high/ba ), .a(\I0/high/latch ), 
        .b(pullcd), .c(\I0/high/latch ), .d(\I0/high/ba ), .e(pullcd), .f(
        \I0/high/ba ) );
    aoi222_1 \I0/high/U1664/U28/U30/U1  ( .x(\I0/high/U1664/x[3] ), .a(
        \I0/high/ncd[7] ), .b(\I0/high/ncd[6] ), .c(\I0/high/ncd[7] ), .d(
        \I0/high/U1664/U28/Z ), .e(\I0/high/ncd[6] ), .f(\I0/high/U1664/U28/Z 
        ) );
    inv_1 \I0/high/U1664/U28/U30/Uinv  ( .x(\I0/high/U1664/U28/Z ), .a(
        \I0/high/U1664/x[3] ) );
    aoi222_1 \I0/high/U1664/U32/U30/U1  ( .x(\I0/high/U1664/x[0] ), .a(
        \I0/high/ncd[1] ), .b(\I0/high/ncd[0] ), .c(\I0/high/ncd[1] ), .d(
        \I0/high/U1664/U32/Z ), .e(\I0/high/ncd[0] ), .f(\I0/high/U1664/U32/Z 
        ) );
    inv_1 \I0/high/U1664/U32/U30/Uinv  ( .x(\I0/high/U1664/U32/Z ), .a(
        \I0/high/U1664/x[0] ) );
    aoi222_1 \I0/high/U1664/U29/U30/U1  ( .x(\I0/high/U1664/x[2] ), .a(
        \I0/high/ncd[5] ), .b(\I0/high/ncd[4] ), .c(\I0/high/ncd[5] ), .d(
        \I0/high/U1664/U29/Z ), .e(\I0/high/ncd[4] ), .f(\I0/high/U1664/U29/Z 
        ) );
    inv_1 \I0/high/U1664/U29/U30/Uinv  ( .x(\I0/high/U1664/U29/Z ), .a(
        \I0/high/U1664/x[2] ) );
    aoi222_1 \I0/high/U1664/U33/U30/U1  ( .x(\I0/high/U1664/y[0] ), .a(
        \I0/high/U1664/x[1] ), .b(\I0/high/U1664/x[0] ), .c(
        \I0/high/U1664/x[1] ), .d(\I0/high/U1664/U33/Z ), .e(
        \I0/high/U1664/x[0] ), .f(\I0/high/U1664/U33/Z ) );
    inv_1 \I0/high/U1664/U33/U30/Uinv  ( .x(\I0/high/U1664/U33/Z ), .a(
        \I0/high/U1664/y[0] ) );
    aoi222_1 \I0/high/U1664/U30/U30/U1  ( .x(\I0/high/U1664/y[1] ), .a(
        \I0/high/U1664/x[3] ), .b(\I0/high/U1664/x[2] ), .c(
        \I0/high/U1664/x[3] ), .d(\I0/high/U1664/U30/Z ), .e(
        \I0/high/U1664/x[2] ), .f(\I0/high/U1664/U30/Z ) );
    inv_1 \I0/high/U1664/U30/U30/Uinv  ( .x(\I0/high/U1664/U30/Z ), .a(
        \I0/high/U1664/y[1] ) );
    aoi222_1 \I0/high/U1664/U31/U30/U1  ( .x(\I0/high/U1664/x[1] ), .a(
        \I0/high/ncd[3] ), .b(\I0/high/ncd[2] ), .c(\I0/high/ncd[3] ), .d(
        \I0/high/U1664/U31/Z ), .e(\I0/high/ncd[2] ), .f(\I0/high/U1664/U31/Z 
        ) );
    inv_1 \I0/high/U1664/U31/U30/Uinv  ( .x(\I0/high/U1664/U31/Z ), .a(
        \I0/high/U1664/x[1] ) );
    aoi222_1 \I0/high/U1664/U37/U30/U1  ( .x(\I0/high/localcd ), .a(
        \I0/high/U1664/y[0] ), .b(\I0/high/U1664/y[1] ), .c(
        \I0/high/U1664/y[0] ), .d(\I0/high/U1664/U37/Z ), .e(
        \I0/high/U1664/y[1] ), .f(\I0/high/U1664/U37/Z ) );
    inv_1 \I0/high/U1664/U37/U30/Uinv  ( .x(\I0/high/U1664/U37/Z ), .a(
        \I0/high/localcd ) );
    nor3_1 \I0/high/U1669/Unr  ( .x(\I0/high/U1669/nr ), .a(
        \I0/high/ctrlack_internal ), .b(n10), .c(\I0/high/drivel ) );
    nand3_1 \I0/high/U1669/Und  ( .x(\I0/high/U1669/nd ), .a(
        \I0/high/ctrlack_internal ), .b(\I0/high/driveh ), .c(\I0/high/drivel 
        ) );
    oa21_1 \I0/high/U1669/U1  ( .x(\I0/high/U1669/n2 ), .a(\I0/high/U1669/n2 ), 
        .b(\I0/high/U1669/nr ), .c(\I0/high/U1669/nd ) );
    inv_2 \I0/high/U1669/U3  ( .x(\I0/net20 ), .a(\I0/high/U1669/n2 ) );
    nor2_1 \I1/U3/U5  ( .x(net31), .a(\I1/net32 ), .b(\I1/net33 ) );
    buf_2 \I1/low/U1653  ( .x(\I1/low/latch ), .a(\I1/net32 ) );
    nor2_1 \I1/low/U264/U5  ( .x(\I1/low/nlocalcd ), .a(reset), .b(
        \I1/low/localcd ) );
    nor2_1 \I1/low/U1659_0_/U5  ( .x(\I1/low/ncd[0] ), .a(ol[16]), .b(oh[16])
         );
    nor2_1 \I1/low/U1659_1_/U5  ( .x(\I1/low/ncd[1] ), .a(ol[17]), .b(oh[17])
         );
    nor2_1 \I1/low/U1659_2_/U5  ( .x(\I1/low/ncd[2] ), .a(ol[18]), .b(oh[18])
         );
    nor2_1 \I1/low/U1659_3_/U5  ( .x(\I1/low/ncd[3] ), .a(ol[19]), .b(oh[19])
         );
    nor2_1 \I1/low/U1659_4_/U5  ( .x(\I1/low/ncd[4] ), .a(ol[20]), .b(oh[20])
         );
    nor2_1 \I1/low/U1659_5_/U5  ( .x(\I1/low/ncd[5] ), .a(ol[21]), .b(oh[21])
         );
    nor2_1 \I1/low/U1659_6_/U5  ( .x(\I1/low/ncd[6] ), .a(ol[22]), .b(oh[22])
         );
    nor2_1 \I1/low/U1659_7_/U5  ( .x(\I1/low/ncd[7] ), .a(ol[23]), .b(oh[23])
         );
    nor2_1 \I1/low/U3/U5  ( .x(\I1/low/ctrlack_internal ), .a(\I1/low/acb ), 
        .b(\I1/low/ba ) );
    buf_2 \I1/low/U1665/U7  ( .x(\I1/low/driveh ), .a(\I1/net20 ) );
    buf_2 \I1/low/U1666/U7  ( .x(\I1/low/drivel ), .a(\I1/net20 ) );
    ao23_1 \I1/low/U1658_0_/U21/U1/U1  ( .x(ol[16]), .a(n8), .b(ol[16]), .c(
        \I1/low/drivel ), .d(pull_l[0]), .e(n7) );
    ao23_1 \I1/low/U1658_1_/U21/U1/U1  ( .x(ol[17]), .a(n8), .b(ol[17]), .c(
        \I1/low/driveh ), .d(pull_l[1]), .e(n7) );
    ao23_1 \I1/low/U1658_2_/U21/U1/U1  ( .x(ol[18]), .a(\I1/low/driveh ), .b(
        ol[18]), .c(n8), .d(pull_l[2]), .e(n7) );
    ao23_1 \I1/low/U1658_3_/U21/U1/U1  ( .x(ol[19]), .a(n8), .b(ol[19]), .c(
        \I1/low/driveh ), .d(pull_l[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_4_/U21/U1/U1  ( .x(ol[20]), .a(\I1/low/drivel ), .b(
        ol[20]), .c(n8), .d(pull_l[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_5_/U21/U1/U1  ( .x(ol[21]), .a(\I1/low/drivel ), .b(
        ol[21]), .c(n8), .d(pull_l[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_6_/U21/U1/U1  ( .x(ol[22]), .a(\I1/low/driveh ), .b(
        ol[22]), .c(\I1/low/drivel ), .d(pull_l[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_7_/U21/U1/U1  ( .x(ol[23]), .a(\I1/low/driveh ), .b(
        ol[23]), .c(\I1/low/driveh ), .d(pull_l[7]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_0_/U21/U1/U1  ( .x(oh[16]), .a(\I1/low/drivel ), .b(
        oh[16]), .c(n8), .d(pull_h[0]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_1_/U21/U1/U1  ( .x(oh[17]), .a(\I1/low/driveh ), .b(
        oh[17]), .c(\I1/low/drivel ), .d(pull_h[1]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_2_/U21/U1/U1  ( .x(oh[18]), .a(\I1/low/drivel ), .b(
        oh[18]), .c(\I1/low/drivel ), .d(pull_h[2]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_3_/U21/U1/U1  ( .x(oh[19]), .a(\I1/low/driveh ), .b(
        oh[19]), .c(\I1/low/driveh ), .d(pull_h[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_4_/U21/U1/U1  ( .x(oh[20]), .a(\I1/low/drivel ), .b(
        oh[20]), .c(\I1/low/driveh ), .d(pull_h[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_5_/U21/U1/U1  ( .x(oh[21]), .a(\I1/low/driveh ), .b(
        oh[21]), .c(n8), .d(pull_h[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_6_/U21/U1/U1  ( .x(oh[22]), .a(n8), .b(oh[22]), .c(
        \I1/low/drivel ), .d(pull_h[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_7_/U21/U1/U1  ( .x(oh[23]), .a(n8), .b(oh[23]), .c(n8
        ), .d(pull_h[7]), .e(\I1/low/latch ) );
    aoai211_1 \I1/low/U4/U28/U1/U1  ( .x(\I1/low/U4/U28/U1/clr ), .a(
        \I1/net20 ), .b(\I1/low/acb ), .c(\I1/low/nlocalcd ), .d(\I1/net32 )
         );
    nand3_1 \I1/low/U4/U28/U1/U2  ( .x(\I1/low/U4/U28/U1/set ), .a(
        \I1/low/nlocalcd ), .b(\I1/net20 ), .c(\I1/low/acb ) );
    nand2_2 \I1/low/U4/U28/U1/U3  ( .x(\I1/net32 ), .a(\I1/low/U4/U28/U1/clr ), 
        .b(\I1/low/U4/U28/U1/set ) );
    oai21_1 \I1/low/U1/U30/U1/U1  ( .x(\I1/low/acb ), .a(\I1/low/U1/Z ), .b(
        \I1/low/ba ), .c(\I1/net20 ) );
    inv_1 \I1/low/U1/U30/U1/U2  ( .x(\I1/low/U1/Z ), .a(\I1/low/acb ) );
    ao222_1 \I1/low/U5/U18/U1/U1  ( .x(\I1/low/ba ), .a(\I1/low/latch ), .b(
        pullcd), .c(\I1/low/latch ), .d(\I1/low/ba ), .e(pullcd), .f(
        \I1/low/ba ) );
    aoi222_1 \I1/low/U1664/U28/U30/U1  ( .x(\I1/low/U1664/x[3] ), .a(
        \I1/low/ncd[7] ), .b(\I1/low/ncd[6] ), .c(\I1/low/ncd[7] ), .d(
        \I1/low/U1664/U28/Z ), .e(\I1/low/ncd[6] ), .f(\I1/low/U1664/U28/Z )
         );
    inv_1 \I1/low/U1664/U28/U30/Uinv  ( .x(\I1/low/U1664/U28/Z ), .a(
        \I1/low/U1664/x[3] ) );
    aoi222_1 \I1/low/U1664/U32/U30/U1  ( .x(\I1/low/U1664/x[0] ), .a(
        \I1/low/ncd[1] ), .b(\I1/low/ncd[0] ), .c(\I1/low/ncd[1] ), .d(
        \I1/low/U1664/U32/Z ), .e(\I1/low/ncd[0] ), .f(\I1/low/U1664/U32/Z )
         );
    inv_1 \I1/low/U1664/U32/U30/Uinv  ( .x(\I1/low/U1664/U32/Z ), .a(
        \I1/low/U1664/x[0] ) );
    aoi222_1 \I1/low/U1664/U29/U30/U1  ( .x(\I1/low/U1664/x[2] ), .a(
        \I1/low/ncd[5] ), .b(\I1/low/ncd[4] ), .c(\I1/low/ncd[5] ), .d(
        \I1/low/U1664/U29/Z ), .e(\I1/low/ncd[4] ), .f(\I1/low/U1664/U29/Z )
         );
    inv_1 \I1/low/U1664/U29/U30/Uinv  ( .x(\I1/low/U1664/U29/Z ), .a(
        \I1/low/U1664/x[2] ) );
    aoi222_1 \I1/low/U1664/U33/U30/U1  ( .x(\I1/low/U1664/y[0] ), .a(
        \I1/low/U1664/x[1] ), .b(\I1/low/U1664/x[0] ), .c(\I1/low/U1664/x[1] ), 
        .d(\I1/low/U1664/U33/Z ), .e(\I1/low/U1664/x[0] ), .f(
        \I1/low/U1664/U33/Z ) );
    inv_1 \I1/low/U1664/U33/U30/Uinv  ( .x(\I1/low/U1664/U33/Z ), .a(
        \I1/low/U1664/y[0] ) );
    aoi222_1 \I1/low/U1664/U30/U30/U1  ( .x(\I1/low/U1664/y[1] ), .a(
        \I1/low/U1664/x[3] ), .b(\I1/low/U1664/x[2] ), .c(\I1/low/U1664/x[3] ), 
        .d(\I1/low/U1664/U30/Z ), .e(\I1/low/U1664/x[2] ), .f(
        \I1/low/U1664/U30/Z ) );
    inv_1 \I1/low/U1664/U30/U30/Uinv  ( .x(\I1/low/U1664/U30/Z ), .a(
        \I1/low/U1664/y[1] ) );
    aoi222_1 \I1/low/U1664/U31/U30/U1  ( .x(\I1/low/U1664/x[1] ), .a(
        \I1/low/ncd[3] ), .b(\I1/low/ncd[2] ), .c(\I1/low/ncd[3] ), .d(
        \I1/low/U1664/U31/Z ), .e(\I1/low/ncd[2] ), .f(\I1/low/U1664/U31/Z )
         );
    inv_1 \I1/low/U1664/U31/U30/Uinv  ( .x(\I1/low/U1664/U31/Z ), .a(
        \I1/low/U1664/x[1] ) );
    aoi222_1 \I1/low/U1664/U37/U30/U1  ( .x(\I1/low/localcd ), .a(
        \I1/low/U1664/y[0] ), .b(\I1/low/U1664/y[1] ), .c(\I1/low/U1664/y[0] ), 
        .d(\I1/low/U1664/U37/Z ), .e(\I1/low/U1664/y[1] ), .f(
        \I1/low/U1664/U37/Z ) );
    inv_1 \I1/low/U1664/U37/U30/Uinv  ( .x(\I1/low/U1664/U37/Z ), .a(
        \I1/low/localcd ) );
    nor3_1 \I1/low/U1669/Unr  ( .x(\I1/low/U1669/nr ), .a(
        \I1/low/ctrlack_internal ), .b(n8), .c(\I1/low/drivel ) );
    nand3_1 \I1/low/U1669/Und  ( .x(\I1/low/U1669/nd ), .a(
        \I1/low/ctrlack_internal ), .b(\I1/low/driveh ), .c(\I1/low/drivel )
         );
    oa21_1 \I1/low/U1669/U1  ( .x(\I1/low/U1669/n2 ), .a(\I1/low/U1669/n2 ), 
        .b(\I1/low/U1669/nr ), .c(\I1/low/U1669/nd ) );
    inv_2 \I1/low/U1669/U3  ( .x(net17), .a(\I1/low/U1669/n2 ) );
    buf_2 \I1/high/U1653  ( .x(\I1/high/latch ), .a(\I1/net33 ) );
    nor2_1 \I1/high/U264/U5  ( .x(\I1/high/nlocalcd ), .a(reset), .b(
        \I1/high/localcd ) );
    nor2_1 \I1/high/U1659_0_/U5  ( .x(\I1/high/ncd[0] ), .a(ol[24]), .b(oh[24]
        ) );
    nor2_1 \I1/high/U1659_1_/U5  ( .x(\I1/high/ncd[1] ), .a(ol[25]), .b(oh[25]
        ) );
    nor2_1 \I1/high/U1659_2_/U5  ( .x(\I1/high/ncd[2] ), .a(ol[26]), .b(oh[26]
        ) );
    nor2_1 \I1/high/U1659_3_/U5  ( .x(\I1/high/ncd[3] ), .a(ol[27]), .b(oh[27]
        ) );
    nor2_1 \I1/high/U1659_4_/U5  ( .x(\I1/high/ncd[4] ), .a(ol[28]), .b(oh[28]
        ) );
    nor2_1 \I1/high/U1659_5_/U5  ( .x(\I1/high/ncd[5] ), .a(ol[29]), .b(oh[29]
        ) );
    nor2_1 \I1/high/U1659_6_/U5  ( .x(\I1/high/ncd[6] ), .a(ol[30]), .b(oh[30]
        ) );
    nor2_1 \I1/high/U1659_7_/U5  ( .x(\I1/high/ncd[7] ), .a(ol[31]), .b(oh[31]
        ) );
    nor2_1 \I1/high/U3/U5  ( .x(\I1/high/ctrlack_internal ), .a(\I1/high/acb ), 
        .b(\I1/high/ba ) );
    ao23_1 \I1/high/U1658_0_/U21/U1/U1  ( .x(ol[24]), .a(n5), .b(ol[24]), .c(
        n6), .d(pull_l[0]), .e(n1) );
    ao23_1 \I1/high/U1658_1_/U21/U1/U1  ( .x(ol[25]), .a(n5), .b(ol[25]), .c(
        n6), .d(pull_l[1]), .e(n1) );
    ao23_1 \I1/high/U1658_2_/U21/U1/U1  ( .x(ol[26]), .a(n5), .b(ol[26]), .c(
        n6), .d(pull_l[2]), .e(n1) );
    ao23_1 \I1/high/U1658_3_/U21/U1/U1  ( .x(ol[27]), .a(n5), .b(ol[27]), .c(
        n5), .d(pull_l[3]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_4_/U21/U1/U1  ( .x(ol[28]), .a(n5), .b(ol[28]), .c(
        n6), .d(pull_l[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_5_/U21/U1/U1  ( .x(ol[29]), .a(n5), .b(ol[29]), .c(
        n6), .d(pull_l[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_6_/U21/U1/U1  ( .x(ol[30]), .a(n5), .b(ol[30]), .c(
        n5), .d(pull_l[6]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_7_/U21/U1/U1  ( .x(ol[31]), .a(n5), .b(ol[31]), .c(
        n5), .d(pull_l[7]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_0_/U21/U1/U1  ( .x(oh[24]), .a(n2), .b(oh[24]), .c(
        n3), .d(pull_h[0]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_1_/U21/U1/U1  ( .x(oh[25]), .a(n2), .b(oh[25]), .c(
        n2), .d(pull_h[1]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_2_/U21/U1/U1  ( .x(oh[26]), .a(n2), .b(oh[26]), .c(
        n3), .d(pull_h[2]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_3_/U21/U1/U1  ( .x(oh[27]), .a(n2), .b(oh[27]), .c(
        n2), .d(pull_h[3]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_4_/U21/U1/U1  ( .x(oh[28]), .a(n2), .b(oh[28]), .c(
        n3), .d(pull_h[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_5_/U21/U1/U1  ( .x(oh[29]), .a(n2), .b(oh[29]), .c(
        n2), .d(pull_h[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_6_/U21/U1/U1  ( .x(oh[30]), .a(n2), .b(oh[30]), .c(
        n3), .d(pull_h[6]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_7_/U21/U1/U1  ( .x(oh[31]), .a(n2), .b(oh[31]), .c(
        n3), .d(pull_h[7]), .e(\I1/high/latch ) );
    aoai211_1 \I1/high/U4/U28/U1/U1  ( .x(\I1/high/U4/U28/U1/clr ), .a(ctrlreq
        ), .b(\I1/high/acb ), .c(\I1/high/nlocalcd ), .d(\I1/net33 ) );
    nand3_1 \I1/high/U4/U28/U1/U2  ( .x(\I1/high/U4/U28/U1/set ), .a(
        \I1/high/nlocalcd ), .b(ctrlreq), .c(\I1/high/acb ) );
    nand2_2 \I1/high/U4/U28/U1/U3  ( .x(\I1/net33 ), .a(
        \I1/high/U4/U28/U1/clr ), .b(\I1/high/U4/U28/U1/set ) );
    oai21_1 \I1/high/U1/U30/U1/U1  ( .x(\I1/high/acb ), .a(\I1/high/U1/Z ), 
        .b(\I1/high/ba ), .c(ctrlreq) );
    inv_1 \I1/high/U1/U30/U1/U2  ( .x(\I1/high/U1/Z ), .a(\I1/high/acb ) );
    ao222_1 \I1/high/U5/U18/U1/U1  ( .x(\I1/high/ba ), .a(\I1/high/latch ), 
        .b(pullcd), .c(\I1/high/latch ), .d(\I1/high/ba ), .e(pullcd), .f(
        \I1/high/ba ) );
    aoi222_1 \I1/high/U1664/U28/U30/U1  ( .x(\I1/high/U1664/x[3] ), .a(
        \I1/high/ncd[7] ), .b(\I1/high/ncd[6] ), .c(\I1/high/ncd[7] ), .d(
        \I1/high/U1664/U28/Z ), .e(\I1/high/ncd[6] ), .f(\I1/high/U1664/U28/Z 
        ) );
    inv_1 \I1/high/U1664/U28/U30/Uinv  ( .x(\I1/high/U1664/U28/Z ), .a(
        \I1/high/U1664/x[3] ) );
    aoi222_1 \I1/high/U1664/U32/U30/U1  ( .x(\I1/high/U1664/x[0] ), .a(
        \I1/high/ncd[1] ), .b(\I1/high/ncd[0] ), .c(\I1/high/ncd[1] ), .d(
        \I1/high/U1664/U32/Z ), .e(\I1/high/ncd[0] ), .f(\I1/high/U1664/U32/Z 
        ) );
    inv_1 \I1/high/U1664/U32/U30/Uinv  ( .x(\I1/high/U1664/U32/Z ), .a(
        \I1/high/U1664/x[0] ) );
    aoi222_1 \I1/high/U1664/U29/U30/U1  ( .x(\I1/high/U1664/x[2] ), .a(
        \I1/high/ncd[5] ), .b(\I1/high/ncd[4] ), .c(\I1/high/ncd[5] ), .d(
        \I1/high/U1664/U29/Z ), .e(\I1/high/ncd[4] ), .f(\I1/high/U1664/U29/Z 
        ) );
    inv_1 \I1/high/U1664/U29/U30/Uinv  ( .x(\I1/high/U1664/U29/Z ), .a(
        \I1/high/U1664/x[2] ) );
    aoi222_1 \I1/high/U1664/U33/U30/U1  ( .x(\I1/high/U1664/y[0] ), .a(
        \I1/high/U1664/x[1] ), .b(\I1/high/U1664/x[0] ), .c(
        \I1/high/U1664/x[1] ), .d(\I1/high/U1664/U33/Z ), .e(
        \I1/high/U1664/x[0] ), .f(\I1/high/U1664/U33/Z ) );
    inv_1 \I1/high/U1664/U33/U30/Uinv  ( .x(\I1/high/U1664/U33/Z ), .a(
        \I1/high/U1664/y[0] ) );
    aoi222_1 \I1/high/U1664/U30/U30/U1  ( .x(\I1/high/U1664/y[1] ), .a(
        \I1/high/U1664/x[3] ), .b(\I1/high/U1664/x[2] ), .c(
        \I1/high/U1664/x[3] ), .d(\I1/high/U1664/U30/Z ), .e(
        \I1/high/U1664/x[2] ), .f(\I1/high/U1664/U30/Z ) );
    inv_1 \I1/high/U1664/U30/U30/Uinv  ( .x(\I1/high/U1664/U30/Z ), .a(
        \I1/high/U1664/y[1] ) );
    aoi222_1 \I1/high/U1664/U31/U30/U1  ( .x(\I1/high/U1664/x[1] ), .a(
        \I1/high/ncd[3] ), .b(\I1/high/ncd[2] ), .c(\I1/high/ncd[3] ), .d(
        \I1/high/U1664/U31/Z ), .e(\I1/high/ncd[2] ), .f(\I1/high/U1664/U31/Z 
        ) );
    inv_1 \I1/high/U1664/U31/U30/Uinv  ( .x(\I1/high/U1664/U31/Z ), .a(
        \I1/high/U1664/x[1] ) );
    aoi222_1 \I1/high/U1664/U37/U30/U1  ( .x(\I1/high/localcd ), .a(
        \I1/high/U1664/y[0] ), .b(\I1/high/U1664/y[1] ), .c(
        \I1/high/U1664/y[0] ), .d(\I1/high/U1664/U37/Z ), .e(
        \I1/high/U1664/y[1] ), .f(\I1/high/U1664/U37/Z ) );
    inv_1 \I1/high/U1664/U37/U30/Uinv  ( .x(\I1/high/U1664/U37/Z ), .a(
        \I1/high/localcd ) );
    nor3_1 \I1/high/U1669/Unr  ( .x(\I1/high/U1669/nr ), .a(
        \I1/high/ctrlack_internal ), .b(n6), .c(n3) );
    nand3_1 \I1/high/U1669/Und  ( .x(\I1/high/U1669/nd ), .a(
        \I1/high/ctrlack_internal ), .b(n6), .c(n3) );
    oa21_1 \I1/high/U1669/U1  ( .x(\I1/high/U1669/n2 ), .a(\I1/high/U1669/n2 ), 
        .b(\I1/high/U1669/nr ), .c(\I1/high/U1669/nd ) );
    inv_2 \I1/high/U1669/U3  ( .x(\I1/net20 ), .a(\I1/high/U1669/n2 ) );
    buf_1 U1 ( .x(n1), .a(\I1/high/latch ) );
    inv_2 U2 ( .x(n2), .a(n4) );
    inv_1 U3 ( .x(n3), .a(n4) );
    inv_0 U4 ( .x(n4), .a(ctrlreq) );
    inv_2 U5 ( .x(n5), .a(n4) );
    inv_1 U6 ( .x(n6), .a(n4) );
    buf_1 U7 ( .x(n7), .a(\I1/low/latch ) );
    buf_2 U8 ( .x(n8), .a(\I1/net20 ) );
    buf_1 U9 ( .x(n9), .a(\I0/high/latch ) );
    buf_2 U10 ( .x(n10), .a(net17) );
    buf_1 U11 ( .x(n11), .a(\I0/low/latch ) );
    buf_2 U12 ( .x(n12), .a(\I0/net20 ) );
endmodule


module chain_fr2dr_byte_0 ( nia, oh, ol, i, nReset, noa );
output [7:0] oh;
output [7:0] ol;
input  [4:0] i;
input  nReset, noa;
output nia;
    wire eop, net135, nca, nbReset, ncla, \c[3] , \c[2] , \c[1] , \c[0] , 
        \cl[3] , \cl[2] , \cl[1] , \cl[0] , asel, bsel, asela, bsela, csel, 
        dsel, csela, dsela, esel, fsel, esela, fsela, naa, nda, \a[3] , \a[2] , 
        \a[1] , \a[0] , \d[3] , \d[2] , \d[1] , \d[0] , nba, nea, nfa, \b[3] , 
        \b[2] , \b[1] , \b[0] , \f[3] , \f[2] , \f[1] , \f[0] , \e[3] , \e[2] , 
        \e[1] , \e[0] , \U891/nack , \U891/acka , \U891/naack[0] , 
        \U891/naack[1] , \U891/iay , \U891/ackb , \U891/reset , \U891/neopack , 
        \U891/U1128/nb , \U891/U1128/na , \U891/U1118_0_/nr , 
        \U891/U1118_0_/nd , \U891/U1118_0_/n2 , \U891/U1118_1_/nr , 
        \U891/U1118_1_/nd , \U891/U1118_1_/n2 , \U891/U1118_2_/nr , 
        \U891/U1118_2_/nd , \U891/U1118_2_/n2 , \U891/U1118_3_/nr , 
        \U891/U1118_3_/nd , \U891/U1118_3_/n2 , \U891/U1117_0_/nr , 
        \U891/U1117_0_/nd , \U891/U1117_0_/n2 , \U891/U1117_1_/nr , 
        \U891/U1117_1_/nd , \U891/U1117_1_/n2 , \U891/U1117_2_/nr , 
        \U891/U1117_2_/nd , \U891/U1117_2_/n2 , \U891/U1117_3_/nr , 
        \U891/U1117_3_/nd , \U891/U1117_3_/n2 , \U886/nack , \U886/acka , 
        \U886/ackb , \U886/reset , \U886/U1128/nb , \U886/U1128/na , 
        \U886/U1127/n5 , \U886/U1127/n1 , \U886/U1127/n2 , \U886/U1127/n3 , 
        \U886/U1127/n4 , \U886/U1118_0_/nr , \U886/U1118_0_/nd , 
        \U886/U1118_0_/n2 , \U886/U1118_1_/nr , \U886/U1118_1_/nd , 
        \U886/U1118_1_/n2 , \U886/U1118_2_/nr , \U886/U1118_2_/nd , 
        \U886/U1118_2_/n2 , \U886/U1118_3_/nr , \U886/U1118_3_/nd , 
        \U886/U1118_3_/n2 , \U886/U1117_0_/nr , \U886/U1117_0_/nd , 
        \U886/U1117_0_/n2 , \U886/U1117_1_/nr , \U886/U1117_1_/nd , 
        \U886/U1117_1_/n2 , \U886/U1117_2_/nr , \U886/U1117_2_/nd , 
        \U886/U1117_2_/n2 , \U886/U1117_3_/nr , \U886/U1117_3_/nd , 
        \U886/U1117_3_/n2 , \U884/nack , \U884/acka , \U884/ackb , 
        \U884/reset , \U884/U1128/nb , \U884/U1128/na , \U884/U1127/n5 , 
        \U884/U1127/n1 , \U884/U1127/n2 , \U884/U1127/n3 , \U884/U1127/n4 , 
        \U884/U1118_0_/nr , \U884/U1118_0_/nd , \U884/U1118_0_/n2 , 
        \U884/U1118_1_/nr , \U884/U1118_1_/nd , \U884/U1118_1_/n2 , 
        \U884/U1118_2_/nr , \U884/U1118_2_/nd , \U884/U1118_2_/n2 , 
        \U884/U1118_3_/nr , \U884/U1118_3_/nd , \U884/U1118_3_/n2 , 
        \U884/U1117_0_/nr , \U884/U1117_0_/nd , \U884/U1117_0_/n2 , 
        \U884/U1117_1_/nr , \U884/U1117_1_/nd , \U884/U1117_1_/n2 , 
        \U884/U1117_2_/nr , \U884/U1117_2_/nd , \U884/U1117_2_/n2 , 
        \U884/U1117_3_/nr , \U884/U1117_3_/nd , \U884/U1117_3_/n2 , 
        \U888/naack , \U888/r , \U888/s , \U888/nback , \U888/reset , 
        \U887/naack , \U887/r , \U887/s , \U887/nback , \U887/reset , 
        \U885/naack , \U885/r , \U885/s , \U885/nback , \U885/reset , \U877/x , 
        \U877/y , \U877/reset , \U877/U590/U25/U1/clr , \U877/U590/U25/U1/ob , 
        \U877/U589/U25/U1/clr , \U877/U589/U25/U1/ob , \U877/U588/U25/U1/clr , 
        \U877/U588/U25/U1/ob , \U877/U591/U25/U1/clr , \U877/U591/U25/U1/ob , 
        \U876/x , \U876/y , \U876/reset , \U876/U590/U25/U1/clr , 
        \U876/U590/U25/U1/ob , \U876/U589/U25/U1/clr , \U876/U589/U25/U1/ob , 
        \U876/U588/U25/U1/clr , \U876/U588/U25/U1/ob , \U876/U591/U25/U1/clr , 
        \U876/U591/U25/U1/ob , \U2/x , \U2/y , \U2/reset , 
        \U2/U590/U25/U1/clr , \U2/U590/U25/U1/ob , \U2/U589/U25/U1/clr , 
        \U2/U589/U25/U1/ob , \U2/U588/U25/U1/clr , \U2/U588/U25/U1/ob , 
        \U2/U591/U25/U1/clr , \U2/U591/U25/U1/ob , \U1/x , \U1/y , \U1/reset , 
        \U1/U590/U25/U1/clr , \U1/U590/U25/U1/ob , \U1/U589/U25/U1/clr , 
        \U1/U589/U25/U1/ob , \U1/U588/U25/U1/clr , \U1/U588/U25/U1/ob , 
        \U1/U591/U25/U1/clr , \U1/U591/U25/U1/ob , \U881/nack[1] , 
        \U881/nack[0] , n1;
    buf_2 U897 ( .x(nbReset), .a(nReset) );
    and4_1 \U894/U12  ( .x(eop), .a(ncla), .b(csela), .c(asela), .d(i[4]) );
    inv_1 \U891/U1126/U3  ( .x(\U891/reset ), .a(nbReset) );
    inv_1 \U891/U1139/U3  ( .x(\U891/neopack ), .a(eop) );
    nand3_1 \U891/U1131/U9  ( .x(\U891/iay ), .a(\U891/neopack ), .b(
        \U891/naack[0] ), .c(\U891/naack[1] ) );
    nor3_1 \U891/U1128/U27  ( .x(\U891/U1128/nb ), .a(\U891/reset ), .b(\b[3] 
        ), .c(\b[2] ) );
    nor2_1 \U891/U1128/U26  ( .x(\U891/U1128/na ), .a(\b[1] ), .b(\b[0] ) );
    nand2_2 \U891/U1128/U29  ( .x(\U891/ackb ), .a(\U891/U1128/nb ), .b(
        \U891/U1128/na ) );
    nor2_1 \U891/U1133/U5  ( .x(\U891/naack[0] ), .a(\a[3] ), .b(\a[2] ) );
    nor2_1 \U891/U1108/U5  ( .x(\U891/nack ), .a(\U891/acka ), .b(\U891/ackb )
         );
    nor2_1 \U891/U1134/U5  ( .x(\U891/naack[1] ), .a(\a[1] ), .b(\a[0] ) );
    nor2_2 \U891/U914/U6  ( .x(nia), .a(\U891/iay ), .b(\U891/ackb ) );
    nand2_1 \U891/U1130/U5  ( .x(\U891/acka ), .a(\U891/naack[0] ), .b(
        \U891/naack[1] ) );
    ao222_4 \U891/U1121/U1/U1  ( .x(bsela), .a(\U891/nack ), .b(bsel), .c(
        \U891/nack ), .d(bsela), .e(bsel), .f(bsela) );
    ao222_4 \U891/U1120/U1/U1  ( .x(asela), .a(asel), .b(\U891/nack ), .c(asel
        ), .d(asela), .e(\U891/nack ), .f(asela) );
    nor3_1 \U891/U1118_0_/Unr  ( .x(\U891/U1118_0_/nr ), .a(i[0]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_0_/Und  ( .x(\U891/U1118_0_/nd ), .a(i[0]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_0_/U1  ( .x(\U891/U1118_0_/n2 ), .a(\U891/U1118_0_/n2 ), 
        .b(\U891/U1118_0_/nr ), .c(\U891/U1118_0_/nd ) );
    inv_2 \U891/U1118_0_/U3  ( .x(\a[0] ), .a(\U891/U1118_0_/n2 ) );
    nor3_1 \U891/U1118_1_/Unr  ( .x(\U891/U1118_1_/nr ), .a(i[1]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_1_/Und  ( .x(\U891/U1118_1_/nd ), .a(i[1]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_1_/U1  ( .x(\U891/U1118_1_/n2 ), .a(\U891/U1118_1_/n2 ), 
        .b(\U891/U1118_1_/nr ), .c(\U891/U1118_1_/nd ) );
    inv_2 \U891/U1118_1_/U3  ( .x(\a[1] ), .a(\U891/U1118_1_/n2 ) );
    nor3_1 \U891/U1118_2_/Unr  ( .x(\U891/U1118_2_/nr ), .a(i[2]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_2_/Und  ( .x(\U891/U1118_2_/nd ), .a(i[2]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_2_/U1  ( .x(\U891/U1118_2_/n2 ), .a(\U891/U1118_2_/n2 ), 
        .b(\U891/U1118_2_/nr ), .c(\U891/U1118_2_/nd ) );
    inv_2 \U891/U1118_2_/U3  ( .x(\a[2] ), .a(\U891/U1118_2_/n2 ) );
    nor3_1 \U891/U1118_3_/Unr  ( .x(\U891/U1118_3_/nr ), .a(i[3]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_3_/Und  ( .x(\U891/U1118_3_/nd ), .a(i[3]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_3_/U1  ( .x(\U891/U1118_3_/n2 ), .a(\U891/U1118_3_/n2 ), 
        .b(\U891/U1118_3_/nr ), .c(\U891/U1118_3_/nd ) );
    inv_2 \U891/U1118_3_/U3  ( .x(\a[3] ), .a(\U891/U1118_3_/n2 ) );
    nor3_1 \U891/U1117_0_/Unr  ( .x(\U891/U1117_0_/nr ), .a(i[0]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_0_/Und  ( .x(\U891/U1117_0_/nd ), .a(i[0]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_0_/U1  ( .x(\U891/U1117_0_/n2 ), .a(\U891/U1117_0_/n2 ), 
        .b(\U891/U1117_0_/nr ), .c(\U891/U1117_0_/nd ) );
    inv_2 \U891/U1117_0_/U3  ( .x(\b[0] ), .a(\U891/U1117_0_/n2 ) );
    nor3_1 \U891/U1117_1_/Unr  ( .x(\U891/U1117_1_/nr ), .a(i[1]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_1_/Und  ( .x(\U891/U1117_1_/nd ), .a(i[1]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_1_/U1  ( .x(\U891/U1117_1_/n2 ), .a(\U891/U1117_1_/n2 ), 
        .b(\U891/U1117_1_/nr ), .c(\U891/U1117_1_/nd ) );
    inv_2 \U891/U1117_1_/U3  ( .x(\b[1] ), .a(\U891/U1117_1_/n2 ) );
    nor3_1 \U891/U1117_2_/Unr  ( .x(\U891/U1117_2_/nr ), .a(i[2]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_2_/Und  ( .x(\U891/U1117_2_/nd ), .a(i[2]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_2_/U1  ( .x(\U891/U1117_2_/n2 ), .a(\U891/U1117_2_/n2 ), 
        .b(\U891/U1117_2_/nr ), .c(\U891/U1117_2_/nd ) );
    inv_2 \U891/U1117_2_/U3  ( .x(\b[2] ), .a(\U891/U1117_2_/n2 ) );
    nor3_1 \U891/U1117_3_/Unr  ( .x(\U891/U1117_3_/nr ), .a(i[3]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_3_/Und  ( .x(\U891/U1117_3_/nd ), .a(i[3]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_3_/U1  ( .x(\U891/U1117_3_/n2 ), .a(\U891/U1117_3_/n2 ), 
        .b(\U891/U1117_3_/nr ), .c(\U891/U1117_3_/nd ) );
    inv_2 \U891/U1117_3_/U3  ( .x(\b[3] ), .a(\U891/U1117_3_/n2 ) );
    inv_1 \U886/U1126/U3  ( .x(\U886/reset ), .a(nbReset) );
    nor3_1 \U886/U1128/U27  ( .x(\U886/U1128/nb ), .a(\U886/reset ), .b(\f[3] 
        ), .c(\f[2] ) );
    nor2_1 \U886/U1128/U26  ( .x(\U886/U1128/na ), .a(\f[1] ), .b(\f[0] ) );
    nand2_2 \U886/U1128/U29  ( .x(\U886/ackb ), .a(\U886/U1128/nb ), .b(
        \U886/U1128/na ) );
    nor2_1 \U886/U1108/U5  ( .x(\U886/nack ), .a(\U886/acka ), .b(\U886/ackb )
         );
    nor2_2 \U886/U914/U6  ( .x(nba), .a(\U886/acka ), .b(\U886/ackb ) );
    and4_1 \U886/U1127/U25  ( .x(\U886/U1127/n5 ), .a(\U886/U1127/n1 ), .b(
        \U886/U1127/n2 ), .c(\U886/U1127/n3 ), .d(\U886/U1127/n4 ) );
    inv_1 \U886/U1127/U1  ( .x(\U886/U1127/n1 ), .a(\e[3] ) );
    inv_1 \U886/U1127/U2  ( .x(\U886/U1127/n2 ), .a(\e[2] ) );
    inv_1 \U886/U1127/U3  ( .x(\U886/U1127/n3 ), .a(\e[1] ) );
    inv_1 \U886/U1127/U4  ( .x(\U886/U1127/n4 ), .a(\e[0] ) );
    inv_2 \U886/U1127/U5  ( .x(\U886/acka ), .a(\U886/U1127/n5 ) );
    ao222_2 \U886/U1121/U19/U1/U1  ( .x(fsela), .a(\U886/nack ), .b(fsel), .c(
        \U886/nack ), .d(fsela), .e(fsel), .f(fsela) );
    ao222_2 \U886/U1120/U19/U1/U1  ( .x(esela), .a(esel), .b(\U886/nack ), .c(
        esel), .d(esela), .e(\U886/nack ), .f(esela) );
    nor3_1 \U886/U1118_0_/Unr  ( .x(\U886/U1118_0_/nr ), .a(\b[0] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_0_/Und  ( .x(\U886/U1118_0_/nd ), .a(\b[0] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_0_/U1  ( .x(\U886/U1118_0_/n2 ), .a(\U886/U1118_0_/n2 ), 
        .b(\U886/U1118_0_/nr ), .c(\U886/U1118_0_/nd ) );
    inv_2 \U886/U1118_0_/U3  ( .x(\e[0] ), .a(\U886/U1118_0_/n2 ) );
    nor3_1 \U886/U1118_1_/Unr  ( .x(\U886/U1118_1_/nr ), .a(\b[1] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_1_/Und  ( .x(\U886/U1118_1_/nd ), .a(\b[1] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_1_/U1  ( .x(\U886/U1118_1_/n2 ), .a(\U886/U1118_1_/n2 ), 
        .b(\U886/U1118_1_/nr ), .c(\U886/U1118_1_/nd ) );
    inv_2 \U886/U1118_1_/U3  ( .x(\e[1] ), .a(\U886/U1118_1_/n2 ) );
    nor3_1 \U886/U1118_2_/Unr  ( .x(\U886/U1118_2_/nr ), .a(\b[2] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_2_/Und  ( .x(\U886/U1118_2_/nd ), .a(\b[2] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_2_/U1  ( .x(\U886/U1118_2_/n2 ), .a(\U886/U1118_2_/n2 ), 
        .b(\U886/U1118_2_/nr ), .c(\U886/U1118_2_/nd ) );
    inv_2 \U886/U1118_2_/U3  ( .x(\e[2] ), .a(\U886/U1118_2_/n2 ) );
    nor3_1 \U886/U1118_3_/Unr  ( .x(\U886/U1118_3_/nr ), .a(\b[3] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_3_/Und  ( .x(\U886/U1118_3_/nd ), .a(\b[3] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_3_/U1  ( .x(\U886/U1118_3_/n2 ), .a(\U886/U1118_3_/n2 ), 
        .b(\U886/U1118_3_/nr ), .c(\U886/U1118_3_/nd ) );
    inv_2 \U886/U1118_3_/U3  ( .x(\e[3] ), .a(\U886/U1118_3_/n2 ) );
    nor3_1 \U886/U1117_0_/Unr  ( .x(\U886/U1117_0_/nr ), .a(\b[0] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_0_/Und  ( .x(\U886/U1117_0_/nd ), .a(\b[0] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_0_/U1  ( .x(\U886/U1117_0_/n2 ), .a(\U886/U1117_0_/n2 ), 
        .b(\U886/U1117_0_/nr ), .c(\U886/U1117_0_/nd ) );
    inv_2 \U886/U1117_0_/U3  ( .x(\f[0] ), .a(\U886/U1117_0_/n2 ) );
    nor3_1 \U886/U1117_1_/Unr  ( .x(\U886/U1117_1_/nr ), .a(\b[1] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_1_/Und  ( .x(\U886/U1117_1_/nd ), .a(\b[1] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_1_/U1  ( .x(\U886/U1117_1_/n2 ), .a(\U886/U1117_1_/n2 ), 
        .b(\U886/U1117_1_/nr ), .c(\U886/U1117_1_/nd ) );
    inv_2 \U886/U1117_1_/U3  ( .x(\f[1] ), .a(\U886/U1117_1_/n2 ) );
    nor3_1 \U886/U1117_2_/Unr  ( .x(\U886/U1117_2_/nr ), .a(\b[2] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_2_/Und  ( .x(\U886/U1117_2_/nd ), .a(\b[2] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_2_/U1  ( .x(\U886/U1117_2_/n2 ), .a(\U886/U1117_2_/n2 ), 
        .b(\U886/U1117_2_/nr ), .c(\U886/U1117_2_/nd ) );
    inv_2 \U886/U1117_2_/U3  ( .x(\f[2] ), .a(\U886/U1117_2_/n2 ) );
    nor3_1 \U886/U1117_3_/Unr  ( .x(\U886/U1117_3_/nr ), .a(\b[3] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_3_/Und  ( .x(\U886/U1117_3_/nd ), .a(\b[3] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_3_/U1  ( .x(\U886/U1117_3_/n2 ), .a(\U886/U1117_3_/n2 ), 
        .b(\U886/U1117_3_/nr ), .c(\U886/U1117_3_/nd ) );
    inv_2 \U886/U1117_3_/U3  ( .x(\f[3] ), .a(\U886/U1117_3_/n2 ) );
    inv_1 \U884/U1126/U3  ( .x(\U884/reset ), .a(nbReset) );
    nor3_1 \U884/U1128/U27  ( .x(\U884/U1128/nb ), .a(\U884/reset ), .b(\d[3] 
        ), .c(\d[2] ) );
    nor2_1 \U884/U1128/U26  ( .x(\U884/U1128/na ), .a(\d[1] ), .b(\d[0] ) );
    nand2_2 \U884/U1128/U29  ( .x(\U884/ackb ), .a(\U884/U1128/nb ), .b(
        \U884/U1128/na ) );
    nor2_1 \U884/U1108/U5  ( .x(\U884/nack ), .a(\U884/acka ), .b(\U884/ackb )
         );
    nor2_2 \U884/U914/U6  ( .x(naa), .a(\U884/acka ), .b(\U884/ackb ) );
    and4_1 \U884/U1127/U25  ( .x(\U884/U1127/n5 ), .a(\U884/U1127/n1 ), .b(
        \U884/U1127/n2 ), .c(\U884/U1127/n3 ), .d(\U884/U1127/n4 ) );
    inv_1 \U884/U1127/U1  ( .x(\U884/U1127/n1 ), .a(\c[3] ) );
    inv_1 \U884/U1127/U2  ( .x(\U884/U1127/n2 ), .a(\c[2] ) );
    inv_1 \U884/U1127/U3  ( .x(\U884/U1127/n3 ), .a(\c[1] ) );
    inv_1 \U884/U1127/U4  ( .x(\U884/U1127/n4 ), .a(\c[0] ) );
    inv_2 \U884/U1127/U5  ( .x(\U884/acka ), .a(\U884/U1127/n5 ) );
    ao222_2 \U884/U1121/U19/U1/U1  ( .x(dsela), .a(\U884/nack ), .b(dsel), .c(
        \U884/nack ), .d(dsela), .e(dsel), .f(dsela) );
    ao222_2 \U884/U1120/U19/U1/U1  ( .x(csela), .a(csel), .b(\U884/nack ), .c(
        csel), .d(csela), .e(\U884/nack ), .f(csela) );
    nor3_1 \U884/U1118_0_/Unr  ( .x(\U884/U1118_0_/nr ), .a(\a[0] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_0_/Und  ( .x(\U884/U1118_0_/nd ), .a(\a[0] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_0_/U1  ( .x(\U884/U1118_0_/n2 ), .a(\U884/U1118_0_/n2 ), 
        .b(\U884/U1118_0_/nr ), .c(\U884/U1118_0_/nd ) );
    inv_2 \U884/U1118_0_/U3  ( .x(\c[0] ), .a(\U884/U1118_0_/n2 ) );
    nor3_1 \U884/U1118_1_/Unr  ( .x(\U884/U1118_1_/nr ), .a(\a[1] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_1_/Und  ( .x(\U884/U1118_1_/nd ), .a(\a[1] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_1_/U1  ( .x(\U884/U1118_1_/n2 ), .a(\U884/U1118_1_/n2 ), 
        .b(\U884/U1118_1_/nr ), .c(\U884/U1118_1_/nd ) );
    inv_2 \U884/U1118_1_/U3  ( .x(\c[1] ), .a(\U884/U1118_1_/n2 ) );
    nor3_1 \U884/U1118_2_/Unr  ( .x(\U884/U1118_2_/nr ), .a(\a[2] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_2_/Und  ( .x(\U884/U1118_2_/nd ), .a(\a[2] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_2_/U1  ( .x(\U884/U1118_2_/n2 ), .a(\U884/U1118_2_/n2 ), 
        .b(\U884/U1118_2_/nr ), .c(\U884/U1118_2_/nd ) );
    inv_2 \U884/U1118_2_/U3  ( .x(\c[2] ), .a(\U884/U1118_2_/n2 ) );
    nor3_1 \U884/U1118_3_/Unr  ( .x(\U884/U1118_3_/nr ), .a(\a[3] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_3_/Und  ( .x(\U884/U1118_3_/nd ), .a(\a[3] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_3_/U1  ( .x(\U884/U1118_3_/n2 ), .a(\U884/U1118_3_/n2 ), 
        .b(\U884/U1118_3_/nr ), .c(\U884/U1118_3_/nd ) );
    inv_2 \U884/U1118_3_/U3  ( .x(\c[3] ), .a(\U884/U1118_3_/n2 ) );
    nor3_1 \U884/U1117_0_/Unr  ( .x(\U884/U1117_0_/nr ), .a(\a[0] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_0_/Und  ( .x(\U884/U1117_0_/nd ), .a(\a[0] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_0_/U1  ( .x(\U884/U1117_0_/n2 ), .a(\U884/U1117_0_/n2 ), 
        .b(\U884/U1117_0_/nr ), .c(\U884/U1117_0_/nd ) );
    inv_2 \U884/U1117_0_/U3  ( .x(\d[0] ), .a(\U884/U1117_0_/n2 ) );
    nor3_1 \U884/U1117_1_/Unr  ( .x(\U884/U1117_1_/nr ), .a(\a[1] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_1_/Und  ( .x(\U884/U1117_1_/nd ), .a(\a[1] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_1_/U1  ( .x(\U884/U1117_1_/n2 ), .a(\U884/U1117_1_/n2 ), 
        .b(\U884/U1117_1_/nr ), .c(\U884/U1117_1_/nd ) );
    inv_2 \U884/U1117_1_/U3  ( .x(\d[1] ), .a(\U884/U1117_1_/n2 ) );
    nor3_1 \U884/U1117_2_/Unr  ( .x(\U884/U1117_2_/nr ), .a(\a[2] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_2_/Und  ( .x(\U884/U1117_2_/nd ), .a(\a[2] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_2_/U1  ( .x(\U884/U1117_2_/n2 ), .a(\U884/U1117_2_/n2 ), 
        .b(\U884/U1117_2_/nr ), .c(\U884/U1117_2_/nd ) );
    inv_2 \U884/U1117_2_/U3  ( .x(\d[2] ), .a(\U884/U1117_2_/n2 ) );
    nor3_1 \U884/U1117_3_/Unr  ( .x(\U884/U1117_3_/nr ), .a(\a[3] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_3_/Und  ( .x(\U884/U1117_3_/nd ), .a(\a[3] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_3_/U1  ( .x(\U884/U1117_3_/n2 ), .a(\U884/U1117_3_/n2 ), 
        .b(\U884/U1117_3_/nr ), .c(\U884/U1117_3_/nd ) );
    inv_2 \U884/U1117_3_/U3  ( .x(\d[3] ), .a(\U884/U1117_3_/n2 ) );
    nand2_1 \U888/U1128/U5  ( .x(\U888/s ), .a(\U888/r ), .b(\U888/nback ) );
    nand2_1 \U888/U1103/U5  ( .x(\U888/r ), .a(\U888/naack ), .b(\U888/s ) );
    inv_1 \U888/U1111/U3  ( .x(\U888/reset ), .a(nbReset) );
    inv_1 \U888/U1112/U3  ( .x(\U888/naack ), .a(esela) );
    nor2_1 \U888/U1127/U5  ( .x(\U888/nback ), .a(fsela), .b(\U888/reset ) );
    and2_2 \U888/U1129/U8  ( .x(esel), .a(\U888/nback ), .b(\U888/s ) );
    and2_2 \U888/U1124/U8  ( .x(fsel), .a(\U888/r ), .b(\U888/naack ) );
    nand2_1 \U887/U1128/U5  ( .x(\U887/s ), .a(\U887/r ), .b(\U887/nback ) );
    nand2_1 \U887/U1103/U5  ( .x(\U887/r ), .a(\U887/naack ), .b(\U887/s ) );
    inv_1 \U887/U1111/U3  ( .x(\U887/reset ), .a(nbReset) );
    inv_1 \U887/U1112/U3  ( .x(\U887/naack ), .a(csela) );
    nor2_1 \U887/U1127/U5  ( .x(\U887/nback ), .a(dsela), .b(\U887/reset ) );
    and2_2 \U887/U1129/U8  ( .x(csel), .a(\U887/nback ), .b(\U887/s ) );
    and2_2 \U887/U1124/U8  ( .x(dsel), .a(\U887/r ), .b(\U887/naack ) );
    nand2_1 \U885/U1128/U5  ( .x(\U885/s ), .a(\U885/r ), .b(\U885/nback ) );
    nand2_1 \U885/U1103/U5  ( .x(\U885/r ), .a(\U885/naack ), .b(\U885/s ) );
    inv_1 \U885/U1111/U3  ( .x(\U885/reset ), .a(nbReset) );
    inv_1 \U885/U1112/U3  ( .x(\U885/naack ), .a(asela) );
    nor2_1 \U885/U1127/U5  ( .x(\U885/nback ), .a(bsela), .b(\U885/reset ) );
    and2_2 \U885/U1129/U8  ( .x(asel), .a(\U885/nback ), .b(\U885/s ) );
    and2_2 \U885/U1124/U8  ( .x(bsel), .a(\U885/r ), .b(\U885/naack ) );
    nor3_1 \U877/U594/U7  ( .x(\U877/x ), .a(ol[7]), .b(\U877/reset ), .c(oh
        [7]) );
    nor3_1 \U877/U593/U7  ( .x(\U877/y ), .a(ol[6]), .b(\U877/reset ), .c(oh
        [6]) );
    inv_1 \U877/U604/U3  ( .x(\U877/reset ), .a(nbReset) );
    oa31_1 \U877/U590/U25/U1/Uclr  ( .x(\U877/U590/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[1] ), .d(oh[6]) );
    oaoi211_1 \U877/U590/U25/U1/Uaoi  ( .x(\U877/U590/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[1] ), .c(n1), .d(\U877/U590/U25/U1/clr ) );
    inv_2 \U877/U590/U25/U1/Ui  ( .x(oh[6]), .a(\U877/U590/U25/U1/ob ) );
    oa31_1 \U877/U589/U25/U1/Uclr  ( .x(\U877/U589/U25/U1/clr ), .a(net135), 
        .b(\cl[1] ), .c(\cl[0] ), .d(ol[7]) );
    oaoi211_1 \U877/U589/U25/U1/Uaoi  ( .x(\U877/U589/U25/U1/ob ), .a(\cl[1] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U589/U25/U1/clr ) );
    inv_2 \U877/U589/U25/U1/Ui  ( .x(ol[7]), .a(\U877/U589/U25/U1/ob ) );
    oa31_1 \U877/U588/U25/U1/Uclr  ( .x(\U877/U588/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[2] ), .d(oh[7]) );
    oaoi211_1 \U877/U588/U25/U1/Uaoi  ( .x(\U877/U588/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[2] ), .c(n1), .d(\U877/U588/U25/U1/clr ) );
    inv_2 \U877/U588/U25/U1/Ui  ( .x(oh[7]), .a(\U877/U588/U25/U1/ob ) );
    oa31_1 \U877/U591/U25/U1/Uclr  ( .x(\U877/U591/U25/U1/clr ), .a(net135), 
        .b(\cl[2] ), .c(\cl[0] ), .d(ol[6]) );
    oaoi211_1 \U877/U591/U25/U1/Uaoi  ( .x(\U877/U591/U25/U1/ob ), .a(\cl[2] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U591/U25/U1/clr ) );
    inv_2 \U877/U591/U25/U1/Ui  ( .x(ol[6]), .a(\U877/U591/U25/U1/ob ) );
    ao222_2 \U877/U592/U19/U1/U1  ( .x(ncla), .a(\U877/x ), .b(\U877/y ), .c(
        \U877/x ), .d(ncla), .e(\U877/y ), .f(ncla) );
    nor3_1 \U876/U594/U7  ( .x(\U876/x ), .a(ol[3]), .b(\U876/reset ), .c(oh
        [3]) );
    nor3_1 \U876/U593/U7  ( .x(\U876/y ), .a(ol[2]), .b(\U876/reset ), .c(oh
        [2]) );
    inv_1 \U876/U604/U3  ( .x(\U876/reset ), .a(nbReset) );
    oa31_1 \U876/U590/U25/U1/Uclr  ( .x(\U876/U590/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[1] ), .d(oh[2]) );
    oaoi211_1 \U876/U590/U25/U1/Uaoi  ( .x(\U876/U590/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[1] ), .c(n1), .d(\U876/U590/U25/U1/clr ) );
    inv_2 \U876/U590/U25/U1/Ui  ( .x(oh[2]), .a(\U876/U590/U25/U1/ob ) );
    oa31_1 \U876/U589/U25/U1/Uclr  ( .x(\U876/U589/U25/U1/clr ), .a(net135), 
        .b(\d[1] ), .c(\d[0] ), .d(ol[3]) );
    oaoi211_1 \U876/U589/U25/U1/Uaoi  ( .x(\U876/U589/U25/U1/ob ), .a(\d[1] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U589/U25/U1/clr ) );
    inv_2 \U876/U589/U25/U1/Ui  ( .x(ol[3]), .a(\U876/U589/U25/U1/ob ) );
    oa31_1 \U876/U588/U25/U1/Uclr  ( .x(\U876/U588/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[2] ), .d(oh[3]) );
    oaoi211_1 \U876/U588/U25/U1/Uaoi  ( .x(\U876/U588/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[2] ), .c(n1), .d(\U876/U588/U25/U1/clr ) );
    inv_2 \U876/U588/U25/U1/Ui  ( .x(oh[3]), .a(\U876/U588/U25/U1/ob ) );
    oa31_1 \U876/U591/U25/U1/Uclr  ( .x(\U876/U591/U25/U1/clr ), .a(net135), 
        .b(\d[2] ), .c(\d[0] ), .d(ol[2]) );
    oaoi211_1 \U876/U591/U25/U1/Uaoi  ( .x(\U876/U591/U25/U1/ob ), .a(\d[2] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U591/U25/U1/clr ) );
    inv_2 \U876/U591/U25/U1/Ui  ( .x(ol[2]), .a(\U876/U591/U25/U1/ob ) );
    ao222_2 \U876/U592/U19/U1/U1  ( .x(nda), .a(\U876/x ), .b(\U876/y ), .c(
        \U876/x ), .d(nda), .e(\U876/y ), .f(nda) );
    nor3_1 \U2/U594/U7  ( .x(\U2/x ), .a(ol[1]), .b(\U2/reset ), .c(oh[1]) );
    nor3_1 \U2/U593/U7  ( .x(\U2/y ), .a(ol[0]), .b(\U2/reset ), .c(oh[0]) );
    inv_1 \U2/U604/U3  ( .x(\U2/reset ), .a(nbReset) );
    oa31_1 \U2/U590/U25/U1/Uclr  ( .x(\U2/U590/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[1] ), .d(oh[0]) );
    oaoi211_1 \U2/U590/U25/U1/Uaoi  ( .x(\U2/U590/U25/U1/ob ), .a(\f[3] ), .b(
        \f[1] ), .c(n1), .d(\U2/U590/U25/U1/clr ) );
    inv_2 \U2/U590/U25/U1/Ui  ( .x(oh[0]), .a(\U2/U590/U25/U1/ob ) );
    oa31_1 \U2/U589/U25/U1/Uclr  ( .x(\U2/U589/U25/U1/clr ), .a(net135), .b(
        \f[1] ), .c(\f[0] ), .d(ol[1]) );
    oaoi211_1 \U2/U589/U25/U1/Uaoi  ( .x(\U2/U589/U25/U1/ob ), .a(\f[1] ), .b(
        \f[0] ), .c(n1), .d(\U2/U589/U25/U1/clr ) );
    inv_2 \U2/U589/U25/U1/Ui  ( .x(ol[1]), .a(\U2/U589/U25/U1/ob ) );
    oa31_1 \U2/U588/U25/U1/Uclr  ( .x(\U2/U588/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[2] ), .d(oh[1]) );
    oaoi211_1 \U2/U588/U25/U1/Uaoi  ( .x(\U2/U588/U25/U1/ob ), .a(\f[3] ), .b(
        \f[2] ), .c(n1), .d(\U2/U588/U25/U1/clr ) );
    inv_2 \U2/U588/U25/U1/Ui  ( .x(oh[1]), .a(\U2/U588/U25/U1/ob ) );
    oa31_1 \U2/U591/U25/U1/Uclr  ( .x(\U2/U591/U25/U1/clr ), .a(net135), .b(
        \f[2] ), .c(\f[0] ), .d(ol[0]) );
    oaoi211_1 \U2/U591/U25/U1/Uaoi  ( .x(\U2/U591/U25/U1/ob ), .a(\f[2] ), .b(
        \f[0] ), .c(n1), .d(\U2/U591/U25/U1/clr ) );
    inv_2 \U2/U591/U25/U1/Ui  ( .x(ol[0]), .a(\U2/U591/U25/U1/ob ) );
    ao222_2 \U2/U592/U19/U1/U1  ( .x(nfa), .a(\U2/x ), .b(\U2/y ), .c(\U2/x ), 
        .d(nfa), .e(\U2/y ), .f(nfa) );
    nor3_1 \U1/U594/U7  ( .x(\U1/x ), .a(ol[5]), .b(\U1/reset ), .c(oh[5]) );
    nor3_1 \U1/U593/U7  ( .x(\U1/y ), .a(ol[4]), .b(\U1/reset ), .c(oh[4]) );
    inv_1 \U1/U604/U3  ( .x(\U1/reset ), .a(nbReset) );
    oa31_1 \U1/U590/U25/U1/Uclr  ( .x(\U1/U590/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[1] ), .d(oh[4]) );
    oaoi211_1 \U1/U590/U25/U1/Uaoi  ( .x(\U1/U590/U25/U1/ob ), .a(\e[3] ), .b(
        \e[1] ), .c(n1), .d(\U1/U590/U25/U1/clr ) );
    inv_2 \U1/U590/U25/U1/Ui  ( .x(oh[4]), .a(\U1/U590/U25/U1/ob ) );
    oa31_1 \U1/U589/U25/U1/Uclr  ( .x(\U1/U589/U25/U1/clr ), .a(net135), .b(
        \e[1] ), .c(\e[0] ), .d(ol[5]) );
    oaoi211_1 \U1/U589/U25/U1/Uaoi  ( .x(\U1/U589/U25/U1/ob ), .a(\e[1] ), .b(
        \e[0] ), .c(n1), .d(\U1/U589/U25/U1/clr ) );
    inv_2 \U1/U589/U25/U1/Ui  ( .x(ol[5]), .a(\U1/U589/U25/U1/ob ) );
    oa31_1 \U1/U588/U25/U1/Uclr  ( .x(\U1/U588/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[2] ), .d(oh[5]) );
    oaoi211_1 \U1/U588/U25/U1/Uaoi  ( .x(\U1/U588/U25/U1/ob ), .a(\e[3] ), .b(
        \e[2] ), .c(n1), .d(\U1/U588/U25/U1/clr ) );
    inv_2 \U1/U588/U25/U1/Ui  ( .x(oh[5]), .a(\U1/U588/U25/U1/ob ) );
    oa31_1 \U1/U591/U25/U1/Uclr  ( .x(\U1/U591/U25/U1/clr ), .a(net135), .b(
        \e[2] ), .c(\e[0] ), .d(ol[4]) );
    oaoi211_1 \U1/U591/U25/U1/Uaoi  ( .x(\U1/U591/U25/U1/ob ), .a(\e[2] ), .b(
        \e[0] ), .c(n1), .d(\U1/U591/U25/U1/clr ) );
    inv_2 \U1/U591/U25/U1/Ui  ( .x(ol[4]), .a(\U1/U591/U25/U1/ob ) );
    ao222_2 \U1/U592/U19/U1/U1  ( .x(nea), .a(\U1/x ), .b(\U1/y ), .c(\U1/x ), 
        .d(nea), .e(\U1/y ), .f(nea) );
    and3_4 \U881/U20/U9  ( .x(nca), .a(\U881/nack[1] ), .b(\U881/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U881/U18/U5  ( .x(\U881/nack[0] ), .a(\cl[3] ), .b(\cl[0] ) );
    nor2_1 \U881/U19/U5  ( .x(\U881/nack[1] ), .a(\cl[1] ), .b(\cl[2] ) );
    ao222_2 \U881/U15_0_/U19/U1/U1  ( .x(\cl[0] ), .a(\c[0] ), .b(ncla), .c(
        \c[0] ), .d(\cl[0] ), .e(ncla), .f(\cl[0] ) );
    ao222_2 \U881/U15_1_/U19/U1/U1  ( .x(\cl[1] ), .a(\c[1] ), .b(ncla), .c(
        \c[1] ), .d(\cl[1] ), .e(ncla), .f(\cl[1] ) );
    ao222_2 \U881/U15_2_/U19/U1/U1  ( .x(\cl[2] ), .a(\c[2] ), .b(ncla), .c(
        \c[2] ), .d(\cl[2] ), .e(ncla), .f(\cl[2] ) );
    ao222_2 \U881/U15_3_/U19/U1/U1  ( .x(\cl[3] ), .a(\c[3] ), .b(ncla), .c(
        \c[3] ), .d(\cl[3] ), .e(ncla), .f(\cl[3] ) );
    and2_5 U1 ( .x(n1), .a(nbReset), .b(noa) );
    and2_3 U2 ( .x(net135), .a(nbReset), .b(noa) );
endmodule


module chain_dr2fr_byte_3 ( eop_ack, ia, o, eop, ih, il, nReset, noa );
output [4:0] o;
input  [7:0] ih;
input  [7:0] il;
input  eop, nReset, noa;
output eop_ack, ia;
    wire eop_pass, nhighack, nlowack, \twobitack[2] , \twobitack[3] , 
        \twobitack[0] , \twobitack[1] , xsel, ysel, nxa, nyla, nbReset, nya, 
        \y[3] , \y[2] , \y[1] , \y[0] , \yl[3] , \yl[2] , \yl[1] , \yl[0] , 
        \cdh[0] , \cdh[1] , \cdl[0] , \cdl[1] , net193, \cdh[2] , \cdh[3] , 
        \cdl[2] , \cdl[3] , net195, bsel, dsel, nba, bg, nda, dg, asel, csel, 
        naa, ag, nca, cg, \d[3] , \d[2] , \d[1] , \d[0] , \b[3] , \b[2] , 
        \b[1] , \b[0] , \x[3] , \x[2] , \x[1] , \x[0] , \c[3] , \c[2] , \c[1] , 
        \c[0] , \a[3] , \a[2] , \a[1] , \a[0] , net194, net199, \U1018/Z , 
        \U1270/net190 , \U1270/net191 , \U1270/net192 , \U1270/net189 , 
        \U1270/U1141/Z , \U1268/net190 , \U1268/net191 , \U1268/net192 , 
        \U1268/net189 , \U1268/U1141/Z , \U1224/nack[0] , \U1224/nack[1] , 
        \U1224/net4 , \U1224/U1125/U28/U1/clr , \U1224/U1125/U28/U1/set , 
        \U1224/U1122/U28/U1/clr , \U1224/U1122/U28/U1/set , 
        \U1224/U916_0_/U25/U1/clr , \U1224/U916_0_/U25/U1/ob , 
        \U1224/U916_1_/U25/U1/clr , \U1224/U916_1_/U25/U1/ob , 
        \U1224/U916_2_/U25/U1/clr , \U1224/U916_2_/U25/U1/ob , 
        \U1224/U916_3_/U25/U1/clr , \U1224/U916_3_/U25/U1/ob , \U1209/nack[0] , 
        \U1209/nack[1] , \U1209/net4 , \U1209/U1125/U28/U1/clr , 
        \U1209/U1125/U28/U1/set , \U1209/U1122/U28/U1/clr , 
        \U1209/U1122/U28/U1/set , \U1209/U916_0_/U25/U1/clr , 
        \U1209/U916_0_/U25/U1/ob , \U1209/U916_1_/U25/U1/clr , 
        \U1209/U916_1_/U25/U1/ob , \U1209/U916_2_/U25/U1/clr , 
        \U1209/U916_2_/U25/U1/ob , \U1209/U916_3_/U25/U1/clr , 
        \U1209/U916_3_/U25/U1/ob , \U1213/nack[0] , \U1213/nack[1] , 
        \U1213/net4 , \U1213/U1125/U28/U1/clr , \U1213/U1125/U28/U1/set , 
        \U1213/U1122/U28/U1/clr , \U1213/U1122/U28/U1/set , 
        \U1213/U916_0_/U25/U1/clr , \U1213/U916_0_/U25/U1/ob , 
        \U1213/U916_1_/U25/U1/clr , \U1213/U916_1_/U25/U1/ob , 
        \U1213/U916_2_/U25/U1/clr , \U1213/U916_2_/U25/U1/ob , 
        \U1213/U916_3_/U25/U1/clr , \U1213/U916_3_/U25/U1/ob , \U1296/ng , 
        \U1296/U1384/Z , \U1296/U1386/U25/U1/clr , \U1296/U1386/U25/U1/ob , 
        \U1298/ng , \U1298/U1384/Z , \U1298/U1386/U25/U1/clr , 
        \U1298/U1386/U25/U1/ob , \U1306/ng , \U1306/U1384/Z , 
        \U1306/U1386/U25/U1/clr , \U1306/U1386/U25/U1/ob , \U1295/ng , 
        \U1295/U1384/Z , \U1295/U1386/U25/U1/clr , \U1295/U1386/U25/U1/ob , 
        \U1297/s , \U1297/nback , \U1297/r , \U1297/naack , \U1297/reset , 
        \U1297/U1128/U28/U1/clr , \U1297/U1128/U28/U1/set , 
        \U1297/U1127/U28/U1/clr , \U1297/U1127/U28/U1/set , \U1300/s , 
        \U1300/nback , \U1300/r , \U1300/naack , \U1300/reset , 
        \U1300/U1128/U28/U1/clr , \U1300/U1128/U28/U1/set , 
        \U1300/U1127/U28/U1/clr , \U1300/U1127/U28/U1/set , \U1289/bnreset , 
        \U1289/U1150/U28/U1/clr , \U1289/U1150/U28/U1/set , 
        \U1289/U1152/U28/U1/clr , \U1289/U1152/U28/U1/set , 
        \U1289/U1149/U28/U1/clr , \U1289/U1149/U28/U1/set , 
        \U1289/U1151/U28/U1/clr , \U1289/U1151/U28/U1/set , 
        \U1289/U1148/net190 , \U1289/U1148/net191 , \U1289/U1148/net192 , 
        \U1289/U1148/net189 , \U1289/U1148/U1141/Z , \U1271/bnreset , 
        \U1271/U1150/U28/U1/clr , \U1271/U1150/U28/U1/set , 
        \U1271/U1152/U28/U1/clr , \U1271/U1152/U28/U1/set , 
        \U1271/U1149/U28/U1/clr , \U1271/U1149/U28/U1/set , 
        \U1271/U1151/U28/U1/clr , \U1271/U1151/U28/U1/set , 
        \U1271/U1148/net190 , \U1271/U1148/net191 , \U1271/U1148/net192 , 
        \U1271/U1148/net189 , \U1271/U1148/U1141/Z , \U1225/naack , \U1225/r , 
        \U1225/s , \U1225/nback , \U1225/reset , \U1308/nack[1] , 
        \U1308/nack[0] ;
    assign o[4] = eop_ack;
    buf_2 U1231 ( .x(nbReset), .a(nReset) );
    and3_1 \U1194/U9  ( .x(eop_pass), .a(nxa), .b(naa), .c(eop) );
    ao222_1 \U1301/U18/U1/U1  ( .x(nlowack), .a(\twobitack[0] ), .b(
        \twobitack[1] ), .c(\twobitack[0] ), .d(nlowack), .e(\twobitack[1] ), 
        .f(nlowack) );
    ao222_1 \U1302/U18/U1/U1  ( .x(nhighack), .a(\twobitack[2] ), .b(
        \twobitack[3] ), .c(\twobitack[2] ), .d(nhighack), .e(\twobitack[3] ), 
        .f(nhighack) );
    aoi222_1 \U1018/U30/U1  ( .x(ia), .a(nhighack), .b(nlowack), .c(nhighack), 
        .d(\U1018/Z ), .e(nlowack), .f(\U1018/Z ) );
    inv_1 \U1018/U30/Uinv  ( .x(\U1018/Z ), .a(ia) );
    ao222_2 \U1038/U19/U1/U1  ( .x(eop_ack), .a(eop_pass), .b(noa), .c(
        eop_pass), .d(eop_ack), .e(noa), .f(eop_ack) );
    inv_1 \U1270/U1147/U3  ( .x(\U1270/net189 ), .a(nbReset) );
    nor2_1 \U1270/U582/U5  ( .x(\U1270/net192 ), .a(il[4]), .b(ih[4]) );
    nor2_1 \U1270/U580/U5  ( .x(\U1270/net191 ), .a(il[5]), .b(ih[5]) );
    nor2_2 \U1270/U1146/U6  ( .x(net199), .a(\U1270/net190 ), .b(
        \U1270/net189 ) );
    aoi222_1 \U1270/U1141/U30/U1  ( .x(\U1270/net190 ), .a(\U1270/net191 ), 
        .b(\U1270/net192 ), .c(\U1270/net191 ), .d(\U1270/U1141/Z ), .e(
        \U1270/net192 ), .f(\U1270/U1141/Z ) );
    inv_1 \U1270/U1141/U30/Uinv  ( .x(\U1270/U1141/Z ), .a(\U1270/net190 ) );
    inv_1 \U1268/U1147/U3  ( .x(\U1268/net189 ), .a(nbReset) );
    nor2_1 \U1268/U582/U5  ( .x(\U1268/net192 ), .a(il[6]), .b(ih[6]) );
    nor2_1 \U1268/U580/U5  ( .x(\U1268/net191 ), .a(il[7]), .b(ih[7]) );
    nor2_2 \U1268/U1146/U6  ( .x(net194), .a(\U1268/net190 ), .b(
        \U1268/net189 ) );
    aoi222_1 \U1268/U1141/U30/U1  ( .x(\U1268/net190 ), .a(\U1268/net191 ), 
        .b(\U1268/net192 ), .c(\U1268/net191 ), .d(\U1268/U1141/Z ), .e(
        \U1268/net192 ), .f(\U1268/U1141/Z ) );
    inv_1 \U1268/U1141/U30/Uinv  ( .x(\U1268/U1141/Z ), .a(\U1268/net190 ) );
    nor2_1 \U1224/U1128/U5  ( .x(\U1224/nack[0] ), .a(\x[3] ), .b(\x[2] ) );
    nor3_1 \U1224/U1127/U7  ( .x(\U1224/nack[1] ), .a(\x[1] ), .b(\U1224/net4 
        ), .c(\x[0] ) );
    inv_1 \U1224/U907/U3  ( .x(\U1224/net4 ), .a(nbReset) );
    aoai211_1 \U1224/U1125/U28/U1/U1  ( .x(\U1224/U1125/U28/U1/clr ), .a(
        \U1224/nack[1] ), .b(\U1224/nack[0] ), .c(asel), .d(naa) );
    nand3_1 \U1224/U1125/U28/U1/U2  ( .x(\U1224/U1125/U28/U1/set ), .a(asel), 
        .b(\U1224/nack[1] ), .c(\U1224/nack[0] ) );
    nand2_2 \U1224/U1125/U28/U1/U3  ( .x(naa), .a(\U1224/U1125/U28/U1/clr ), 
        .b(\U1224/U1125/U28/U1/set ) );
    aoai211_1 \U1224/U1122/U28/U1/U1  ( .x(\U1224/U1122/U28/U1/clr ), .a(
        \U1224/nack[0] ), .b(\U1224/nack[1] ), .c(csel), .d(nca) );
    nand3_1 \U1224/U1122/U28/U1/U2  ( .x(\U1224/U1122/U28/U1/set ), .a(csel), 
        .b(\U1224/nack[0] ), .c(\U1224/nack[1] ) );
    nand2_2 \U1224/U1122/U28/U1/U3  ( .x(nca), .a(\U1224/U1122/U28/U1/clr ), 
        .b(\U1224/U1122/U28/U1/set ) );
    oa31_1 \U1224/U916_0_/U25/U1/Uclr  ( .x(\U1224/U916_0_/U25/U1/clr ), .a(
        nxa), .b(\a[0] ), .c(\c[0] ), .d(\x[0] ) );
    oaoi211_1 \U1224/U916_0_/U25/U1/Uaoi  ( .x(\U1224/U916_0_/U25/U1/ob ), .a(
        \a[0] ), .b(\c[0] ), .c(nxa), .d(\U1224/U916_0_/U25/U1/clr ) );
    inv_2 \U1224/U916_0_/U25/U1/Ui  ( .x(\x[0] ), .a(\U1224/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_1_/U25/U1/Uclr  ( .x(\U1224/U916_1_/U25/U1/clr ), .a(
        nxa), .b(\a[1] ), .c(\c[1] ), .d(\x[1] ) );
    oaoi211_1 \U1224/U916_1_/U25/U1/Uaoi  ( .x(\U1224/U916_1_/U25/U1/ob ), .a(
        \a[1] ), .b(\c[1] ), .c(nxa), .d(\U1224/U916_1_/U25/U1/clr ) );
    inv_2 \U1224/U916_1_/U25/U1/Ui  ( .x(\x[1] ), .a(\U1224/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_2_/U25/U1/Uclr  ( .x(\U1224/U916_2_/U25/U1/clr ), .a(
        nxa), .b(\a[2] ), .c(\c[2] ), .d(\x[2] ) );
    oaoi211_1 \U1224/U916_2_/U25/U1/Uaoi  ( .x(\U1224/U916_2_/U25/U1/ob ), .a(
        \a[2] ), .b(\c[2] ), .c(nxa), .d(\U1224/U916_2_/U25/U1/clr ) );
    inv_2 \U1224/U916_2_/U25/U1/Ui  ( .x(\x[2] ), .a(\U1224/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_3_/U25/U1/Uclr  ( .x(\U1224/U916_3_/U25/U1/clr ), .a(
        nxa), .b(\a[3] ), .c(\c[3] ), .d(\x[3] ) );
    oaoi211_1 \U1224/U916_3_/U25/U1/Uaoi  ( .x(\U1224/U916_3_/U25/U1/ob ), .a(
        \a[3] ), .b(\c[3] ), .c(nxa), .d(\U1224/U916_3_/U25/U1/clr ) );
    inv_2 \U1224/U916_3_/U25/U1/Ui  ( .x(\x[3] ), .a(\U1224/U916_3_/U25/U1/ob 
        ) );
    nor2_1 \U1209/U1128/U5  ( .x(\U1209/nack[0] ), .a(o[3]), .b(o[2]) );
    nor3_1 \U1209/U1127/U7  ( .x(\U1209/nack[1] ), .a(o[1]), .b(\U1209/net4 ), 
        .c(o[0]) );
    inv_1 \U1209/U907/U3  ( .x(\U1209/net4 ), .a(nbReset) );
    aoai211_1 \U1209/U1125/U28/U1/U1  ( .x(\U1209/U1125/U28/U1/clr ), .a(
        \U1209/nack[1] ), .b(\U1209/nack[0] ), .c(xsel), .d(nxa) );
    nand3_1 \U1209/U1125/U28/U1/U2  ( .x(\U1209/U1125/U28/U1/set ), .a(xsel), 
        .b(\U1209/nack[1] ), .c(\U1209/nack[0] ) );
    nand2_2 \U1209/U1125/U28/U1/U3  ( .x(nxa), .a(\U1209/U1125/U28/U1/clr ), 
        .b(\U1209/U1125/U28/U1/set ) );
    aoai211_1 \U1209/U1122/U28/U1/U1  ( .x(\U1209/U1122/U28/U1/clr ), .a(
        \U1209/nack[0] ), .b(\U1209/nack[1] ), .c(ysel), .d(nyla) );
    nand3_1 \U1209/U1122/U28/U1/U2  ( .x(\U1209/U1122/U28/U1/set ), .a(ysel), 
        .b(\U1209/nack[0] ), .c(\U1209/nack[1] ) );
    nand2_2 \U1209/U1122/U28/U1/U3  ( .x(nyla), .a(\U1209/U1122/U28/U1/clr ), 
        .b(\U1209/U1122/U28/U1/set ) );
    oa31_1 \U1209/U916_0_/U25/U1/Uclr  ( .x(\U1209/U916_0_/U25/U1/clr ), .a(
        noa), .b(\x[0] ), .c(\yl[0] ), .d(o[0]) );
    oaoi211_1 \U1209/U916_0_/U25/U1/Uaoi  ( .x(\U1209/U916_0_/U25/U1/ob ), .a(
        \x[0] ), .b(\yl[0] ), .c(noa), .d(\U1209/U916_0_/U25/U1/clr ) );
    inv_2 \U1209/U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U1209/U916_0_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_1_/U25/U1/Uclr  ( .x(\U1209/U916_1_/U25/U1/clr ), .a(
        noa), .b(\x[1] ), .c(\yl[1] ), .d(o[1]) );
    oaoi211_1 \U1209/U916_1_/U25/U1/Uaoi  ( .x(\U1209/U916_1_/U25/U1/ob ), .a(
        \x[1] ), .b(\yl[1] ), .c(noa), .d(\U1209/U916_1_/U25/U1/clr ) );
    inv_2 \U1209/U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U1209/U916_1_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_2_/U25/U1/Uclr  ( .x(\U1209/U916_2_/U25/U1/clr ), .a(
        noa), .b(\x[2] ), .c(\yl[2] ), .d(o[2]) );
    oaoi211_1 \U1209/U916_2_/U25/U1/Uaoi  ( .x(\U1209/U916_2_/U25/U1/ob ), .a(
        \x[2] ), .b(\yl[2] ), .c(noa), .d(\U1209/U916_2_/U25/U1/clr ) );
    inv_2 \U1209/U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U1209/U916_2_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_3_/U25/U1/Uclr  ( .x(\U1209/U916_3_/U25/U1/clr ), .a(
        noa), .b(\x[3] ), .c(\yl[3] ), .d(o[3]) );
    oaoi211_1 \U1209/U916_3_/U25/U1/Uaoi  ( .x(\U1209/U916_3_/U25/U1/ob ), .a(
        \x[3] ), .b(\yl[3] ), .c(noa), .d(\U1209/U916_3_/U25/U1/clr ) );
    inv_2 \U1209/U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U1209/U916_3_/U25/U1/ob )
         );
    nor2_1 \U1213/U1128/U5  ( .x(\U1213/nack[0] ), .a(\y[3] ), .b(\y[2] ) );
    nor3_1 \U1213/U1127/U7  ( .x(\U1213/nack[1] ), .a(\y[1] ), .b(\U1213/net4 
        ), .c(\y[0] ) );
    inv_1 \U1213/U907/U3  ( .x(\U1213/net4 ), .a(nbReset) );
    aoai211_1 \U1213/U1125/U28/U1/U1  ( .x(\U1213/U1125/U28/U1/clr ), .a(
        \U1213/nack[1] ), .b(\U1213/nack[0] ), .c(bsel), .d(nba) );
    nand3_1 \U1213/U1125/U28/U1/U2  ( .x(\U1213/U1125/U28/U1/set ), .a(bsel), 
        .b(\U1213/nack[1] ), .c(\U1213/nack[0] ) );
    nand2_2 \U1213/U1125/U28/U1/U3  ( .x(nba), .a(\U1213/U1125/U28/U1/clr ), 
        .b(\U1213/U1125/U28/U1/set ) );
    aoai211_1 \U1213/U1122/U28/U1/U1  ( .x(\U1213/U1122/U28/U1/clr ), .a(
        \U1213/nack[0] ), .b(\U1213/nack[1] ), .c(dsel), .d(nda) );
    nand3_1 \U1213/U1122/U28/U1/U2  ( .x(\U1213/U1122/U28/U1/set ), .a(dsel), 
        .b(\U1213/nack[0] ), .c(\U1213/nack[1] ) );
    nand2_2 \U1213/U1122/U28/U1/U3  ( .x(nda), .a(\U1213/U1122/U28/U1/clr ), 
        .b(\U1213/U1122/U28/U1/set ) );
    oa31_1 \U1213/U916_0_/U25/U1/Uclr  ( .x(\U1213/U916_0_/U25/U1/clr ), .a(
        nya), .b(\b[0] ), .c(\d[0] ), .d(\y[0] ) );
    oaoi211_1 \U1213/U916_0_/U25/U1/Uaoi  ( .x(\U1213/U916_0_/U25/U1/ob ), .a(
        \b[0] ), .b(\d[0] ), .c(nya), .d(\U1213/U916_0_/U25/U1/clr ) );
    inv_2 \U1213/U916_0_/U25/U1/Ui  ( .x(\y[0] ), .a(\U1213/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_1_/U25/U1/Uclr  ( .x(\U1213/U916_1_/U25/U1/clr ), .a(
        nya), .b(\b[1] ), .c(\d[1] ), .d(\y[1] ) );
    oaoi211_1 \U1213/U916_1_/U25/U1/Uaoi  ( .x(\U1213/U916_1_/U25/U1/ob ), .a(
        \b[1] ), .b(\d[1] ), .c(nya), .d(\U1213/U916_1_/U25/U1/clr ) );
    inv_2 \U1213/U916_1_/U25/U1/Ui  ( .x(\y[1] ), .a(\U1213/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_2_/U25/U1/Uclr  ( .x(\U1213/U916_2_/U25/U1/clr ), .a(
        nya), .b(\b[2] ), .c(\d[2] ), .d(\y[2] ) );
    oaoi211_1 \U1213/U916_2_/U25/U1/Uaoi  ( .x(\U1213/U916_2_/U25/U1/ob ), .a(
        \b[2] ), .b(\d[2] ), .c(nya), .d(\U1213/U916_2_/U25/U1/clr ) );
    inv_2 \U1213/U916_2_/U25/U1/Ui  ( .x(\y[2] ), .a(\U1213/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_3_/U25/U1/Uclr  ( .x(\U1213/U916_3_/U25/U1/clr ), .a(
        nya), .b(\b[3] ), .c(\d[3] ), .d(\y[3] ) );
    oaoi211_1 \U1213/U916_3_/U25/U1/Uaoi  ( .x(\U1213/U916_3_/U25/U1/ob ), .a(
        \b[3] ), .b(\d[3] ), .c(nya), .d(\U1213/U916_3_/U25/U1/clr ) );
    inv_2 \U1213/U916_3_/U25/U1/Ui  ( .x(\y[3] ), .a(\U1213/U916_3_/U25/U1/ob 
        ) );
    and3_2 \U1210/U1138/U9  ( .x(\d[3] ), .a(\cdh[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1137/U9  ( .x(\d[2] ), .a(\cdl[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1139/U9  ( .x(\d[1] ), .a(\cdh[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1210/U1136/U9  ( .x(\d[0] ), .a(\cdl[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1162/U1138/U9  ( .x(\a[3] ), .a(ih[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1137/U9  ( .x(\a[2] ), .a(il[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1139/U9  ( .x(\a[1] ), .a(ih[6]), .b(naa), .c(il[7]) );
    and3_2 \U1162/U1136/U9  ( .x(\a[0] ), .a(il[6]), .b(naa), .c(il[7]) );
    and3_2 \U1211/U1138/U9  ( .x(\b[3] ), .a(ih[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1137/U9  ( .x(\b[2] ), .a(il[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1139/U9  ( .x(\b[1] ), .a(ih[4]), .b(nba), .c(il[5]) );
    and3_2 \U1211/U1136/U9  ( .x(\b[0] ), .a(il[4]), .b(nba), .c(il[5]) );
    and3_2 \U1163/U1138/U9  ( .x(\c[3] ), .a(\cdh[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1137/U9  ( .x(\c[2] ), .a(\cdl[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1139/U9  ( .x(\c[1] ), .a(\cdh[2] ), .b(nca), .c(\cdl[3] )
         );
    and3_2 \U1163/U1136/U9  ( .x(\c[0] ), .a(\cdl[2] ), .b(nca), .c(\cdl[3] )
         );
    and2_1 \U1296/U1385/U8  ( .x(cg), .a(nbReset), .b(\U1296/ng ) );
    aoi222_1 \U1296/U1384/U30/U1  ( .x(\U1296/ng ), .a(nca), .b(net195), .c(
        nca), .d(\U1296/U1384/Z ), .e(net195), .f(\U1296/U1384/Z ) );
    inv_1 \U1296/U1384/U30/Uinv  ( .x(\U1296/U1384/Z ), .a(\U1296/ng ) );
    oa31_1 \U1296/U1386/U25/U1/Uclr  ( .x(\U1296/U1386/U25/U1/clr ), .a(
        \twobitack[2] ), .b(cg), .c(nca), .d(net195) );
    oaoi211_1 \U1296/U1386/U25/U1/Uaoi  ( .x(\U1296/U1386/U25/U1/ob ), .a(cg), 
        .b(nca), .c(\twobitack[2] ), .d(\U1296/U1386/U25/U1/clr ) );
    inv_2 \U1296/U1386/U25/U1/Ui  ( .x(net195), .a(\U1296/U1386/U25/U1/ob ) );
    and2_1 \U1298/U1385/U8  ( .x(dg), .a(nbReset), .b(\U1298/ng ) );
    aoi222_1 \U1298/U1384/U30/U1  ( .x(\U1298/ng ), .a(nda), .b(net193), .c(
        nda), .d(\U1298/U1384/Z ), .e(net193), .f(\U1298/U1384/Z ) );
    inv_1 \U1298/U1384/U30/Uinv  ( .x(\U1298/U1384/Z ), .a(\U1298/ng ) );
    oa31_1 \U1298/U1386/U25/U1/Uclr  ( .x(\U1298/U1386/U25/U1/clr ), .a(
        \twobitack[0] ), .b(dg), .c(nda), .d(net193) );
    oaoi211_1 \U1298/U1386/U25/U1/Uaoi  ( .x(\U1298/U1386/U25/U1/ob ), .a(dg), 
        .b(nda), .c(\twobitack[0] ), .d(\U1298/U1386/U25/U1/clr ) );
    inv_2 \U1298/U1386/U25/U1/Ui  ( .x(net193), .a(\U1298/U1386/U25/U1/ob ) );
    and2_1 \U1306/U1385/U8  ( .x(bg), .a(nbReset), .b(\U1306/ng ) );
    aoi222_1 \U1306/U1384/U30/U1  ( .x(\U1306/ng ), .a(nba), .b(\twobitack[1] 
        ), .c(nba), .d(\U1306/U1384/Z ), .e(\twobitack[1] ), .f(
        \U1306/U1384/Z ) );
    inv_1 \U1306/U1384/U30/Uinv  ( .x(\U1306/U1384/Z ), .a(\U1306/ng ) );
    oa31_1 \U1306/U1386/U25/U1/Uclr  ( .x(\U1306/U1386/U25/U1/clr ), .a(net199
        ), .b(bg), .c(nba), .d(\twobitack[1] ) );
    oaoi211_1 \U1306/U1386/U25/U1/Uaoi  ( .x(\U1306/U1386/U25/U1/ob ), .a(bg), 
        .b(nba), .c(net199), .d(\U1306/U1386/U25/U1/clr ) );
    inv_2 \U1306/U1386/U25/U1/Ui  ( .x(\twobitack[1] ), .a(
        \U1306/U1386/U25/U1/ob ) );
    and2_1 \U1295/U1385/U8  ( .x(ag), .a(nbReset), .b(\U1295/ng ) );
    aoi222_1 \U1295/U1384/U30/U1  ( .x(\U1295/ng ), .a(naa), .b(\twobitack[3] 
        ), .c(naa), .d(\U1295/U1384/Z ), .e(\twobitack[3] ), .f(
        \U1295/U1384/Z ) );
    inv_1 \U1295/U1384/U30/Uinv  ( .x(\U1295/U1384/Z ), .a(\U1295/ng ) );
    oa31_1 \U1295/U1386/U25/U1/Uclr  ( .x(\U1295/U1386/U25/U1/clr ), .a(net194
        ), .b(ag), .c(naa), .d(\twobitack[3] ) );
    oaoi211_1 \U1295/U1386/U25/U1/Uaoi  ( .x(\U1295/U1386/U25/U1/ob ), .a(ag), 
        .b(naa), .c(net194), .d(\U1295/U1386/U25/U1/clr ) );
    inv_2 \U1295/U1386/U25/U1/Ui  ( .x(\twobitack[3] ), .a(
        \U1295/U1386/U25/U1/ob ) );
    nand2_1 \U1297/U1131/U5  ( .x(\U1297/s ), .a(\U1297/r ), .b(\U1297/nback )
         );
    nand2_1 \U1297/U1103/U5  ( .x(\U1297/r ), .a(\U1297/naack ), .b(\U1297/s )
         );
    inv_1 \U1297/U1111/U3  ( .x(\U1297/reset ), .a(nbReset) );
    inv_1 \U1297/U1112/U3  ( .x(\U1297/naack ), .a(naa) );
    nor2_1 \U1297/U1130/U5  ( .x(\U1297/nback ), .a(nca), .b(\U1297/reset ) );
    aoai211_1 \U1297/U1128/U28/U1/U1  ( .x(\U1297/U1128/U28/U1/clr ), .a(
        \U1297/r ), .b(\U1297/naack ), .c(cg), .d(csel) );
    nand3_1 \U1297/U1128/U28/U1/U2  ( .x(\U1297/U1128/U28/U1/set ), .a(cg), 
        .b(\U1297/r ), .c(\U1297/naack ) );
    nand2_2 \U1297/U1128/U28/U1/U3  ( .x(csel), .a(\U1297/U1128/U28/U1/clr ), 
        .b(\U1297/U1128/U28/U1/set ) );
    aoai211_1 \U1297/U1127/U28/U1/U1  ( .x(\U1297/U1127/U28/U1/clr ), .a(
        \U1297/s ), .b(\U1297/nback ), .c(ag), .d(asel) );
    nand3_1 \U1297/U1127/U28/U1/U2  ( .x(\U1297/U1127/U28/U1/set ), .a(ag), 
        .b(\U1297/s ), .c(\U1297/nback ) );
    nand2_2 \U1297/U1127/U28/U1/U3  ( .x(asel), .a(\U1297/U1127/U28/U1/clr ), 
        .b(\U1297/U1127/U28/U1/set ) );
    nand2_1 \U1300/U1131/U5  ( .x(\U1300/s ), .a(\U1300/r ), .b(\U1300/nback )
         );
    nand2_1 \U1300/U1103/U5  ( .x(\U1300/r ), .a(\U1300/naack ), .b(\U1300/s )
         );
    inv_1 \U1300/U1111/U3  ( .x(\U1300/reset ), .a(nbReset) );
    inv_1 \U1300/U1112/U3  ( .x(\U1300/naack ), .a(nba) );
    nor2_1 \U1300/U1130/U5  ( .x(\U1300/nback ), .a(nda), .b(\U1300/reset ) );
    aoai211_1 \U1300/U1128/U28/U1/U1  ( .x(\U1300/U1128/U28/U1/clr ), .a(
        \U1300/r ), .b(\U1300/naack ), .c(dg), .d(dsel) );
    nand3_1 \U1300/U1128/U28/U1/U2  ( .x(\U1300/U1128/U28/U1/set ), .a(dg), 
        .b(\U1300/r ), .c(\U1300/naack ) );
    nand2_2 \U1300/U1128/U28/U1/U3  ( .x(dsel), .a(\U1300/U1128/U28/U1/clr ), 
        .b(\U1300/U1128/U28/U1/set ) );
    aoai211_1 \U1300/U1127/U28/U1/U1  ( .x(\U1300/U1127/U28/U1/clr ), .a(
        \U1300/s ), .b(\U1300/nback ), .c(bg), .d(bsel) );
    nand3_1 \U1300/U1127/U28/U1/U2  ( .x(\U1300/U1127/U28/U1/set ), .a(bg), 
        .b(\U1300/s ), .c(\U1300/nback ) );
    nand2_2 \U1300/U1127/U28/U1/U3  ( .x(bsel), .a(\U1300/U1127/U28/U1/clr ), 
        .b(\U1300/U1127/U28/U1/set ) );
    aoai211_1 \U1289/U1150/U28/U1/U1  ( .x(\U1289/U1150/U28/U1/clr ), .a(il[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[2] ) );
    nand3_1 \U1289/U1150/U28/U1/U2  ( .x(\U1289/U1150/U28/U1/set ), .a(net195), 
        .b(il[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1150/U28/U1/U3  ( .x(\cdl[2] ), .a(
        \U1289/U1150/U28/U1/clr ), .b(\U1289/U1150/U28/U1/set ) );
    aoai211_1 \U1289/U1152/U28/U1/U1  ( .x(\U1289/U1152/U28/U1/clr ), .a(il[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[3] ) );
    nand3_1 \U1289/U1152/U28/U1/U2  ( .x(\U1289/U1152/U28/U1/set ), .a(net195), 
        .b(il[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1152/U28/U1/U3  ( .x(\cdl[3] ), .a(
        \U1289/U1152/U28/U1/clr ), .b(\U1289/U1152/U28/U1/set ) );
    aoai211_1 \U1289/U1149/U28/U1/U1  ( .x(\U1289/U1149/U28/U1/clr ), .a(ih[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[2] ) );
    nand3_1 \U1289/U1149/U28/U1/U2  ( .x(\U1289/U1149/U28/U1/set ), .a(net195), 
        .b(ih[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1149/U28/U1/U3  ( .x(\cdh[2] ), .a(
        \U1289/U1149/U28/U1/clr ), .b(\U1289/U1149/U28/U1/set ) );
    aoai211_1 \U1289/U1151/U28/U1/U1  ( .x(\U1289/U1151/U28/U1/clr ), .a(ih[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[3] ) );
    nand3_1 \U1289/U1151/U28/U1/U2  ( .x(\U1289/U1151/U28/U1/set ), .a(net195), 
        .b(ih[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1151/U28/U1/U3  ( .x(\cdh[3] ), .a(
        \U1289/U1151/U28/U1/clr ), .b(\U1289/U1151/U28/U1/set ) );
    inv_1 \U1289/U1148/U1147/U3  ( .x(\U1289/U1148/net189 ), .a(
        \U1289/bnreset ) );
    nor2_1 \U1289/U1148/U582/U5  ( .x(\U1289/U1148/net192 ), .a(\cdl[3] ), .b(
        \cdh[3] ) );
    nor2_1 \U1289/U1148/U580/U5  ( .x(\U1289/U1148/net191 ), .a(\cdl[2] ), .b(
        \cdh[2] ) );
    nor2_2 \U1289/U1148/U1146/U6  ( .x(\twobitack[2] ), .a(
        \U1289/U1148/net190 ), .b(\U1289/U1148/net189 ) );
    aoi222_1 \U1289/U1148/U1141/U30/U1  ( .x(\U1289/U1148/net190 ), .a(
        \U1289/U1148/net191 ), .b(\U1289/U1148/net192 ), .c(
        \U1289/U1148/net191 ), .d(\U1289/U1148/U1141/Z ), .e(
        \U1289/U1148/net192 ), .f(\U1289/U1148/U1141/Z ) );
    inv_1 \U1289/U1148/U1141/U30/Uinv  ( .x(\U1289/U1148/U1141/Z ), .a(
        \U1289/U1148/net190 ) );
    aoai211_1 \U1271/U1150/U28/U1/U1  ( .x(\U1271/U1150/U28/U1/clr ), .a(il[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[0] ) );
    nand3_1 \U1271/U1150/U28/U1/U2  ( .x(\U1271/U1150/U28/U1/set ), .a(net193), 
        .b(il[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1150/U28/U1/U3  ( .x(\cdl[0] ), .a(
        \U1271/U1150/U28/U1/clr ), .b(\U1271/U1150/U28/U1/set ) );
    aoai211_1 \U1271/U1152/U28/U1/U1  ( .x(\U1271/U1152/U28/U1/clr ), .a(il[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[1] ) );
    nand3_1 \U1271/U1152/U28/U1/U2  ( .x(\U1271/U1152/U28/U1/set ), .a(net193), 
        .b(il[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1152/U28/U1/U3  ( .x(\cdl[1] ), .a(
        \U1271/U1152/U28/U1/clr ), .b(\U1271/U1152/U28/U1/set ) );
    aoai211_1 \U1271/U1149/U28/U1/U1  ( .x(\U1271/U1149/U28/U1/clr ), .a(ih[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[0] ) );
    nand3_1 \U1271/U1149/U28/U1/U2  ( .x(\U1271/U1149/U28/U1/set ), .a(net193), 
        .b(ih[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1149/U28/U1/U3  ( .x(\cdh[0] ), .a(
        \U1271/U1149/U28/U1/clr ), .b(\U1271/U1149/U28/U1/set ) );
    aoai211_1 \U1271/U1151/U28/U1/U1  ( .x(\U1271/U1151/U28/U1/clr ), .a(ih[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[1] ) );
    nand3_1 \U1271/U1151/U28/U1/U2  ( .x(\U1271/U1151/U28/U1/set ), .a(net193), 
        .b(ih[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1151/U28/U1/U3  ( .x(\cdh[1] ), .a(
        \U1271/U1151/U28/U1/clr ), .b(\U1271/U1151/U28/U1/set ) );
    inv_1 \U1271/U1148/U1147/U3  ( .x(\U1271/U1148/net189 ), .a(
        \U1271/bnreset ) );
    nor2_1 \U1271/U1148/U582/U5  ( .x(\U1271/U1148/net192 ), .a(\cdl[1] ), .b(
        \cdh[1] ) );
    nor2_1 \U1271/U1148/U580/U5  ( .x(\U1271/U1148/net191 ), .a(\cdl[0] ), .b(
        \cdh[0] ) );
    nor2_2 \U1271/U1148/U1146/U6  ( .x(\twobitack[0] ), .a(
        \U1271/U1148/net190 ), .b(\U1271/U1148/net189 ) );
    aoi222_1 \U1271/U1148/U1141/U30/U1  ( .x(\U1271/U1148/net190 ), .a(
        \U1271/U1148/net191 ), .b(\U1271/U1148/net192 ), .c(
        \U1271/U1148/net191 ), .d(\U1271/U1148/U1141/Z ), .e(
        \U1271/U1148/net192 ), .f(\U1271/U1148/U1141/Z ) );
    inv_1 \U1271/U1148/U1141/U30/Uinv  ( .x(\U1271/U1148/U1141/Z ), .a(
        \U1271/U1148/net190 ) );
    nand2_1 \U1225/U1128/U5  ( .x(\U1225/s ), .a(\U1225/r ), .b(\U1225/nback )
         );
    nand2_1 \U1225/U1103/U5  ( .x(\U1225/r ), .a(\U1225/naack ), .b(\U1225/s )
         );
    inv_1 \U1225/U1111/U3  ( .x(\U1225/reset ), .a(nbReset) );
    inv_1 \U1225/U1112/U3  ( .x(\U1225/naack ), .a(nxa) );
    nor2_1 \U1225/U1127/U5  ( .x(\U1225/nback ), .a(nyla), .b(\U1225/reset )
         );
    and2_2 \U1225/U1129/U8  ( .x(xsel), .a(\U1225/nback ), .b(\U1225/s ) );
    and2_2 \U1225/U1124/U8  ( .x(ysel), .a(\U1225/r ), .b(\U1225/naack ) );
    and3_4 \U1308/U20/U9  ( .x(nya), .a(\U1308/nack[1] ), .b(\U1308/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U1308/U18/U5  ( .x(\U1308/nack[0] ), .a(\yl[3] ), .b(\yl[0] ) );
    nor2_1 \U1308/U19/U5  ( .x(\U1308/nack[1] ), .a(\yl[1] ), .b(\yl[2] ) );
    ao222_2 \U1308/U15_0_/U19/U1/U1  ( .x(\yl[0] ), .a(\y[0] ), .b(nyla), .c(
        \y[0] ), .d(\yl[0] ), .e(nyla), .f(\yl[0] ) );
    ao222_2 \U1308/U15_1_/U19/U1/U1  ( .x(\yl[1] ), .a(\y[1] ), .b(nyla), .c(
        \y[1] ), .d(\yl[1] ), .e(nyla), .f(\yl[1] ) );
    ao222_2 \U1308/U15_2_/U19/U1/U1  ( .x(\yl[2] ), .a(\y[2] ), .b(nyla), .c(
        \y[2] ), .d(\yl[2] ), .e(nyla), .f(\yl[2] ) );
    ao222_2 \U1308/U15_3_/U19/U1/U1  ( .x(\yl[3] ), .a(\y[3] ), .b(nyla), .c(
        \y[3] ), .d(\yl[3] ), .e(nyla), .f(\yl[3] ) );
    buf_3 U1 ( .x(\U1271/bnreset ), .a(nbReset) );
    buf_3 U2 ( .x(\U1289/bnreset ), .a(nbReset) );
endmodule


module chain_dr8bit_completion_12 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_13 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_14 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_15 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr32bit_completion_8 ( o, i );
input  [63:0] i;
output o;
    wire nx, \cd[3] , \cd[2] , ny, \cd[0] , \cd[1] , \U16/Z , \U6/Z , \U15/Z ;
    chain_dr8bit_completion_12 U11 ( .o(\cd[3] ), .i({i[63], i[62], i[61], 
        i[60], i[59], i[58], i[57], i[56], i[31], i[30], i[29], i[28], i[27], 
        i[26], i[25], i[24]}) );
    chain_dr8bit_completion_15 U14 ( .o(\cd[2] ), .i({i[55], i[54], i[53], 
        i[52], i[51], i[50], i[49], i[48], i[23], i[22], i[21], i[20], i[19], 
        i[18], i[17], i[16]}) );
    chain_dr8bit_completion_14 U13 ( .o(\cd[1] ), .i({i[47], i[46], i[45], 
        i[44], i[43], i[42], i[41], i[40], i[15], i[14], i[13], i[12], i[11], 
        i[10], i[9], i[8]}) );
    chain_dr8bit_completion_13 U12 ( .o(\cd[0] ), .i({i[39], i[38], i[37], 
        i[36], i[35], i[34], i[33], i[32], i[7], i[6], i[5], i[4], i[3], i[2], 
        i[1], i[0]}) );
    aoi222_1 \U16/U30/U1  ( .x(ny), .a(\cd[0] ), .b(\cd[1] ), .c(\cd[0] ), .d(
        \U16/Z ), .e(\cd[1] ), .f(\U16/Z ) );
    inv_1 \U16/U30/Uinv  ( .x(\U16/Z ), .a(ny) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(ny), .b(nx), .c(ny), .d(\U6/Z ), .e(nx), 
        .f(\U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U15/U30/U1  ( .x(nx), .a(\cd[3] ), .b(\cd[2] ), .c(\cd[3] ), .d(
        \U15/Z ), .e(\cd[2] ), .f(\U15/Z ) );
    inv_1 \U15/U30/Uinv  ( .x(\U15/Z ), .a(nx) );
endmodule


module chain_selement_ga_68 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_69 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_t_ctrl_0 ( cack, fcdefer, fcslowack, screq, ack, defer, fcack, 
    nReset, scack, slowack );
input  ack, defer, fcack, nReset, scack, slowack;
output cack, fcdefer, fcslowack, screq;
    wire net269, net280, net275, net270, net265, net278, net276, net277, 
        net263, net271, net266, net279, net272, net264, net267, net273, net268, 
        net274, \U49/U28/U1/clr , \U49/U28/U1/set , \U50/U28/U1/clr , 
        \U50/U28/U1/set , \U51/U28/U1/clr , \U51/U28/U1/set , \U57/acb , 
        \U57/U1/Z ;
    chain_selement_ga_69 U55 ( .Aa(net269), .Br(fcdefer), .Ar(net280), .Ba(
        fcack) );
    chain_selement_ga_68 U54 ( .Aa(net275), .Br(fcslowack), .Ar(net270), .Ba(
        fcack) );
    or2_4 \U12/U12  ( .x(net268), .a(net266), .b(net270) );
    or2_4 \U56/U12  ( .x(net274), .a(net275), .b(net269) );
    or2_4 \U14/U12  ( .x(net273), .a(net274), .b(net266) );
    or3_1 \U36/U12  ( .x(cack), .a(net267), .b(net264), .c(net272) );
    nor3_1 \U21/U7  ( .x(net271), .a(net270), .b(net266), .c(net280) );
    and2_1 \U53/U8  ( .x(net263), .a(net271), .b(nReset) );
    and2_1 \U43/U8  ( .x(net277), .a(net265), .b(nReset) );
    nor2_1 \U22/U5  ( .x(net265), .a(net278), .b(net276) );
    ao222_2 \U44/U19/U1/U1  ( .x(net276), .a(net280), .b(net273), .c(net280), 
        .d(net276), .e(net273), .f(net276) );
    ao222_2 \U40/U19/U1/U1  ( .x(net280), .a(net272), .b(net277), .c(net272), 
        .d(net280), .e(net277), .f(net280) );
    ao222_2 \U45/U19/U1/U1  ( .x(net279), .a(net273), .b(net268), .c(net273), 
        .d(net279), .e(net268), .f(net279) );
    ao222_2 \U42/U19/U1/U1  ( .x(net266), .a(net277), .b(net267), .c(net277), 
        .d(net266), .e(net267), .f(net266) );
    ao222_2 \U39/U19/U1/U1  ( .x(net270), .a(net277), .b(net264), .c(net277), 
        .d(net270), .e(net264), .f(net270) );
    aoai211_1 \U49/U28/U1/U1  ( .x(\U49/U28/U1/clr ), .a(ack), .b(nReset), .c(
        net263), .d(net267) );
    nand3_1 \U49/U28/U1/U2  ( .x(\U49/U28/U1/set ), .a(net263), .b(ack), .c(
        nReset) );
    nand2_2 \U49/U28/U1/U3  ( .x(net267), .a(\U49/U28/U1/clr ), .b(
        \U49/U28/U1/set ) );
    aoai211_1 \U50/U28/U1/U1  ( .x(\U50/U28/U1/clr ), .a(slowack), .b(nReset), 
        .c(net263), .d(net264) );
    nand3_1 \U50/U28/U1/U2  ( .x(\U50/U28/U1/set ), .a(net263), .b(slowack), 
        .c(nReset) );
    nand2_2 \U50/U28/U1/U3  ( .x(net264), .a(\U50/U28/U1/clr ), .b(
        \U50/U28/U1/set ) );
    aoai211_1 \U51/U28/U1/U1  ( .x(\U51/U28/U1/clr ), .a(defer), .b(nReset), 
        .c(net263), .d(net272) );
    nand2_2 \U51/U28/U1/U3  ( .x(net272), .a(\U51/U28/U1/clr ), .b(
        \U51/U28/U1/set ) );
    and2_1 \U57/U2/U8  ( .x(screq), .a(net279), .b(\U57/acb ) );
    nor2_1 \U57/U3/U5  ( .x(net278), .a(\U57/acb ), .b(scack) );
    oai21_1 \U57/U1/U30/U1/U1  ( .x(\U57/acb ), .a(\U57/U1/Z ), .b(scack), .c(
        net279) );
    inv_1 \U57/U1/U30/U1/U2  ( .x(\U57/U1/Z ), .a(\U57/acb ) );
    nand3_0 U1 ( .x(\U51/U28/U1/set ), .a(net263), .b(defer), .c(nReset) );
endmodule


module chain_mergepackets_3 ( naa, nba, o, a, b, nReset, noa );
output [4:0] o;
input  [4:0] a;
input  [4:0] b;
input  nReset, noa;
output naa, nba;
    wire \noack[1] , \noack[0] , reset, bsel, as, setb, asel, seta, 
        \U916_0_/U25/U1/clr , \U916_0_/U25/U1/ob , \U916_1_/U25/U1/clr , 
        \U916_1_/U25/U1/ob , \U916_2_/U25/U1/clr , \U916_2_/U25/U1/ob , 
        \U916_3_/U25/U1/clr , \U916_3_/U25/U1/ob ;
    and2_1 \U1155/U8  ( .x(as), .a(seta), .b(asel) );
    nand2_1 \U1145/U5  ( .x(asel), .a(bsel), .b(seta) );
    nand2_1 \U1103/U5  ( .x(bsel), .a(setb), .b(asel) );
    inv_1 \U1135/U3  ( .x(reset), .a(nReset) );
    inv_1 \U1134/U3  ( .x(setb), .a(a[4]) );
    and3_2 \U1154/U9  ( .x(naa), .a(\noack[1] ), .b(\noack[0] ), .c(as) );
    nor3_1 \U1127/U7  ( .x(\noack[0] ), .a(o[1]), .b(reset), .c(o[0]) );
    nor2_1 \U1132/U5  ( .x(\noack[1] ), .a(o[3]), .b(o[2]) );
    oa31_1 \U916_0_/U25/U1/Uclr  ( .x(\U916_0_/U25/U1/clr ), .a(noa), .b(a[0]), 
        .c(b[0]), .d(o[0]) );
    oaoi211_1 \U916_0_/U25/U1/Uaoi  ( .x(\U916_0_/U25/U1/ob ), .a(a[0]), .b(b
        [0]), .c(noa), .d(\U916_0_/U25/U1/clr ) );
    inv_2 \U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U916_0_/U25/U1/ob ) );
    oa31_1 \U916_1_/U25/U1/Uclr  ( .x(\U916_1_/U25/U1/clr ), .a(noa), .b(a[1]), 
        .c(b[1]), .d(o[1]) );
    oaoi211_1 \U916_1_/U25/U1/Uaoi  ( .x(\U916_1_/U25/U1/ob ), .a(a[1]), .b(b
        [1]), .c(noa), .d(\U916_1_/U25/U1/clr ) );
    inv_2 \U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U916_1_/U25/U1/ob ) );
    oa31_1 \U916_2_/U25/U1/Uclr  ( .x(\U916_2_/U25/U1/clr ), .a(noa), .b(a[2]), 
        .c(b[2]), .d(o[2]) );
    oaoi211_1 \U916_2_/U25/U1/Uaoi  ( .x(\U916_2_/U25/U1/ob ), .a(a[2]), .b(b
        [2]), .c(noa), .d(\U916_2_/U25/U1/clr ) );
    inv_2 \U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U916_2_/U25/U1/ob ) );
    oa31_1 \U916_3_/U25/U1/Uclr  ( .x(\U916_3_/U25/U1/clr ), .a(noa), .b(a[3]), 
        .c(b[3]), .d(o[3]) );
    oaoi211_1 \U916_3_/U25/U1/Uaoi  ( .x(\U916_3_/U25/U1/ob ), .a(a[3]), .b(b
        [3]), .c(noa), .d(\U916_3_/U25/U1/clr ) );
    inv_2 \U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U916_3_/U25/U1/ob ) );
    ao222_2 \U1148/U19/U1/U1  ( .x(o[4]), .a(noa), .b(b[4]), .c(noa), .d(o[4]), 
        .e(b[4]), .f(o[4]) );
    aoi21_1 \U1153/U11  ( .x(seta), .a(o[4]), .b(setb), .c(reset) );
    and3_3 U1 ( .x(nba), .a(bsel), .b(\noack[0] ), .c(\noack[1] ) );
endmodule


module target_wb ( addr, ccol, chainresponse, crnw, csize, ctag, lock, 
    nchaincommandack, nrouteack, pred, rack, routetxreq, seq, tag_h, tag_l, wd, 
    cack, cdefer, chaincommand, cndefer, cok, err, nReset, nchainresponseack, 
    rd, route, routetxack );
output [63:0] addr;
output [5:0] ccol;
output [4:0] chainresponse;
output [1:0] crnw;
output [3:0] csize;
output [9:0] ctag;
output [1:0] lock;
output [1:0] pred;
output [1:0] seq;
output [4:0] tag_h;
output [4:0] tag_l;
output [63:0] wd;
input  [4:0] chaincommand;
input  [1:0] err;
input  [63:0] rd;
input  [4:0] route;
input  cack, cdefer, cndefer, cok, nReset, nchainresponseack, routetxack;
output nchaincommandack, nrouteack, rack, routetxreq;
    wire n11, n12, n13, n14, n15, \net242[0] , \net242[1] , \net242[2] , 
        \net242[3] , \net242[4] , \net242[5] , \net242[6] , \net242[7] , 
        \net242[8] , \net242[9] , \net242[10] , \net243[0] , \net243[1] , 
        \net243[2] , \net243[3] , \net243[4] , \net243[5] , \net243[6] , 
        \net243[7] , \net243[8] , \net243[9] , \net243[10] , \net244[0] , 
        \net244[1] , \net244[2] , \net244[3] , \net244[4] , \net244[5] , 
        \net244[6] , \net244[7] , \net244[8] , \net244[9] , \net244[10] , 
        \chainff_l[7] , \chainff_l[6] , \chainff_l[5] , \chainff_l[4] , 
        \chainff_l[3] , \chainff_l[2] , \chainff_l[1] , \chainff_l[0] , 
        \chdrack[0] , \chdrack[1] , \obl[7] , \obl[6] , \obl[5] , \obl[4] , 
        \obl[3] , \obl[2] , \obl[1] , \obl[0] , \tcbh[7] , \tcbh[6] , 
        \tcbh[5] , \tcbh[4] , \tcbh[3] , \tcbh[2] , \tcbh[1] , \tcbh[0] , 
        \tcbl[7] , \tcbl[6] , \tcbl[5] , \tcbl[4] , \tcbl[3] , \tcbl[2] , 
        \tcbl[1] , \tcbl[0] , \tresponse[4] , \tresponse[3] , \tresponse[2] , 
        \tresponse[1] , \tresponse[0] , \nchdr_ack[10] , \nchdr_ack[9] , 
        \nchdr_ack[8] , \nchdr_ack[7] , \nchdr_ack[6] , \nchdr_ack[5] , 
        \nchdr_ack[4] , \nchdr_ack[3] , \nchdr_ack[2] , \nchdr_ack[1] , 
        \nchdr_ack[0] , \chainff_h[7] , \chainff_h[6] , \chainff_h[5] , 
        \chainff_h[4] , \chainff_h[3] , \chainff_h[2] , \chainff_h[1] , 
        \chainff_h[0] , \rhdr_l[15] , \rhdr_l[14] , \rhdr_l[13] , \rhdr_l[7] , 
        \rhdr_l[6] , \rhdr_l[5] , \obh[7] , \obh[6] , \obh[5] , \obh[4] , 
        \obh[3] , \obh[2] , \obh[1] , \obh[0] , \rhdr_h[15] , \rhdr_h[14] , 
        \rhdr_h[13] , \rhdr_h[7] , \rhdr_h[6] , \rhdr_h[5] , net265, nbreset, 
        net248, rhdrack, read_ctrlack, chainff_ack, read_req, read_cd, teop, 
        fcack, tcba, net145, screq, fcslowack, fcdefer, read_ack, 
        ntresponseack, net200, noba, pullcd, net168, net188, net201, net194, 
        net178, net189, net191, net284, hdrcd, chdrctrlack, \U1770/U21/nr , 
        \U1770/U21/nd , \U1770/U21/n2 , \U1761/U28/Z , \U1761/U32/Z , 
        \U1761/U29/Z , \U1761/U33/Z , \U1761/U30/Z , \U1761/U31/Z , \U1632/Z , 
        \U1676/Z , \U1761/y[0] , \U1761/y[1] , \U1761/x[1] , \U1761/x[3] , 
        \U1761/x[2] , \U1761/x[0] , \U1574_0_/net231 , \U1574_1_/net231 , 
        \U1574_2_/net231 , \U1574_3_/net231 , \U1574_4_/net231 , 
        \U1574_5_/net231 , \U1574_6_/net231 , \U1574_7_/net231 , 
        \U1574_8_/net231 , \U1574_9_/net231 , \U1574_10_/net231 , n4, n7, n8, 
        n9, n10;
    chain_sendword_0 U1765 ( .ctrlack(read_ctrlack), .oh({\chainff_h[7] , 
        \chainff_h[6] , \chainff_h[5] , \chainff_h[4] , \chainff_h[3] , 
        \chainff_h[2] , \chainff_h[1] , \chainff_h[0] }), .ol({\chainff_l[7] , 
        \chainff_l[6] , \chainff_l[5] , \chainff_l[4] , \chainff_l[3] , 
        \chainff_l[2] , \chainff_l[1] , \chainff_l[0] }), .chainackff(
        chainff_ack), .ctrlreq(read_req), .ih(rd[63:32]), .il(rd[31:0]) );
    chain_dr32bit_completion_8 rd_cd ( .o(read_cd), .i(rd) );
    chain_trhdr_0 xmitHdr ( .chainff_ack(chainff_ack), .chainh({\tcbh[7] , 
        \tcbh[6] , \tcbh[5] , \tcbh[4] , \tcbh[3] , \tcbh[2] , \tcbh[1] , 
        \tcbh[0] }), .chainl({\tcbl[7] , \tcbl[6] , \tcbl[5] , \tcbl[4] , 
        \tcbl[3] , \tcbl[2] , \tcbl[1] , \tcbl[0] }), .eop(teop), .hdrack(
        rhdrack), .normal_ack(rack), .notify_ack(fcack), .read_req(read_req), 
        .routereq(routetxreq), .chain_ff_h({\chainff_h[7] , \chainff_h[6] , 
        \chainff_h[5] , \chainff_h[4] , \chainff_h[3] , \chainff_h[2] , 
        \chainff_h[1] , \chainff_h[0] }), .chainack(tcba), .chainff_l({
        \chainff_l[7] , \chainff_l[6] , \chainff_l[5] , \chainff_l[4] , 
        \chainff_l[3] , \chainff_l[2] , \chainff_l[1] , \chainff_l[0] }), 
        .eopack(net145), .err(err), .nReset(n7), .normal_response(screq), 
        .notify_accept(fcslowack), .notify_defer(fcdefer), .rcol_h({
        \rhdr_h[15] , \rhdr_h[14] , \rhdr_h[13] }), .rcol_l({\rhdr_l[15] , 
        \rhdr_l[14] , \rhdr_l[13] }), .read_ack(read_ack), .rnw_h(\rhdr_h[7] ), 
        .rnw_l(\rhdr_l[7] ), .routeack(routetxack), .rsize_h({\rhdr_h[6] , 
        \rhdr_h[5] }), .rsize_l({\rhdr_l[6] , \rhdr_l[5] }), .rtag_h(tag_h), 
        .rtag_l(tag_l) );
    chain_dr2fr_byte_3 dr2fr ( .eop_ack(net145), .ia(tcba), .o({\tresponse[4] , 
        \tresponse[3] , \tresponse[2] , \tresponse[1] , \tresponse[0] }), 
        .eop(teop), .ih({\tcbh[7] , \tcbh[6] , \tcbh[5] , \tcbh[4] , \tcbh[3] , 
        \tcbh[2] , \tcbh[1] , \tcbh[0] }), .il({\tcbl[7] , \tcbl[6] , 
        \tcbl[5] , \tcbl[4] , \tcbl[3] , \tcbl[2] , \tcbl[1] , \tcbl[0] }), 
        .nReset(nbreset), .noa(ntresponseack) );
    chain_mergepackets_3 merger ( .naa(nrouteack), .nba(ntresponseack), .o(
        chainresponse), .a(route), .b({\tresponse[4] , \tresponse[3] , 
        \tresponse[2] , \tresponse[1] , \tresponse[0] }), .nReset(nbreset), 
        .noa(nchainresponseack) );
    chain_tchdr_0 header ( .addr_req(net200), .col_h(ccol[5:3]), .col_l(ccol
        [2:0]), .itag_h(ctag[9:5]), .itag_l(ctag[4:0]), .lock(lock), .ncback(
        noba), .pred(pred), .pullcd(pullcd), .reset(net168), .rnw_h(n11), 
        .rnw_l(n12), .seq(seq), .size_h({n13, csize[2]}), .size_l({n14, n15}), 
        .write_req(net188), .chwh({\obh[7] , \obh[6] , \obh[5] , \obh[4] , 
        \obh[3] , \obh[2] , \obh[1] , \obh[0] }), .chwl({\obl[7] , \obl[6] , 
        \obl[5] , \obl[4] , \obl[3] , \obl[2] , \obl[1] , \obl[0] }), 
        .addr_ack(net201), .addr_pull(net194), .nReset(n7), .nack(net178), 
        .write_ack(net189), .write_pull(net191) );
    chain_irdemux_32new_1 wd_hld ( .ctrlack(net189), .oh(wd[63:32]), .ol(wd
        [31:0]), .pullreq(net191), .pull_h({\obh[7] , \obh[6] , \obh[5] , 
        \obh[4] , \obh[3] , \obh[2] , \obh[1] , \obh[0] }), .pull_l({\obl[7] , 
        \obl[6] , \obl[5] , \obl[4] , \obl[3] , \obl[2] , \obl[1] , \obl[0] }), 
        .pullcd(pullcd), .reset(net168), .ctrlreq(net188) );
    chain_irdemux_32new_0 adr_hld ( .ctrlack(net201), .oh(addr[63:32]), .ol(
        addr[31:0]), .pullreq(net194), .pull_h({\obh[7] , \obh[6] , \obh[5] , 
        \obh[4] , \obh[3] , \obh[2] , \obh[1] , \obh[0] }), .pull_l({\obl[7] , 
        \obl[6] , \obl[5] , \obl[4] , \obl[3] , \obl[2] , \obl[1] , \obl[0] }), 
        .pullcd(pullcd), .reset(net168), .ctrlreq(net200) );
    chain_fr2dr_byte_0 chain_decoder ( .nia(nchaincommandack), .oh({\obh[7] , 
        \obh[6] , \obh[5] , \obh[4] , \obh[3] , \obh[2] , \obh[1] , \obh[0] }), 
        .ol({\obl[7] , \obl[6] , \obl[5] , \obl[4] , \obl[3] , \obl[2] , 
        \obl[1] , \obl[0] }), .i(chaincommand), .nReset(nbreset), .noa(noba)
         );
    chain_t_ctrl_0 cmd_ctrl ( .cack(net284), .fcdefer(fcdefer), .fcslowack(
        fcslowack), .screq(screq), .ack(cok), .defer(cdefer), .fcack(fcack), 
        .nReset(n7), .scack(rack), .slowack(cndefer) );
    inv_1 \I4/U3  ( .x(net265), .a(nbreset) );
    ao222_1 \U1761/U37/U18/U1/U1  ( .x(\chdrack[0] ), .a(\U1761/y[0] ), .b(
        \U1761/y[1] ), .c(\U1761/y[0] ), .d(\chdrack[0] ), .e(\U1761/y[1] ), 
        .f(\chdrack[0] ) );
    ao222_1 \U1762/U18/U1/U1  ( .x(chdrctrlack), .a(hdrcd), .b(net284), .c(
        hdrcd), .d(chdrctrlack), .e(net284), .f(chdrctrlack) );
    ao222_1 \U1769/U18/U1/U1  ( .x(read_ack), .a(read_ctrlack), .b(read_cd), 
        .c(read_ctrlack), .d(read_ack), .e(read_cd), .f(read_ack) );
    aoi222_1 \U1761/U28/U30/U1  ( .x(\U1761/x[3] ), .a(\nchdr_ack[7] ), .b(
        \nchdr_ack[6] ), .c(\nchdr_ack[7] ), .d(\U1761/U28/Z ), .e(
        \nchdr_ack[6] ), .f(\U1761/U28/Z ) );
    inv_1 \U1761/U28/U30/Uinv  ( .x(\U1761/U28/Z ), .a(\U1761/x[3] ) );
    aoi222_1 \U1761/U32/U30/U1  ( .x(\U1761/x[0] ), .a(\nchdr_ack[1] ), .b(
        \nchdr_ack[0] ), .c(\nchdr_ack[1] ), .d(\U1761/U32/Z ), .e(
        \nchdr_ack[0] ), .f(\U1761/U32/Z ) );
    inv_1 \U1761/U32/U30/Uinv  ( .x(\U1761/U32/Z ), .a(\U1761/x[0] ) );
    aoi222_1 \U1761/U29/U30/U1  ( .x(\U1761/x[2] ), .a(\nchdr_ack[5] ), .b(
        \nchdr_ack[4] ), .c(\nchdr_ack[5] ), .d(\U1761/U29/Z ), .e(
        \nchdr_ack[4] ), .f(\U1761/U29/Z ) );
    inv_1 \U1761/U29/U30/Uinv  ( .x(\U1761/U29/Z ), .a(\U1761/x[2] ) );
    aoi222_1 \U1761/U33/U30/U1  ( .x(\U1761/y[0] ), .a(\U1761/x[1] ), .b(
        \U1761/x[0] ), .c(\U1761/x[1] ), .d(\U1761/U33/Z ), .e(\U1761/x[0] ), 
        .f(\U1761/U33/Z ) );
    inv_1 \U1761/U33/U30/Uinv  ( .x(\U1761/U33/Z ), .a(\U1761/y[0] ) );
    aoi222_1 \U1761/U30/U30/U1  ( .x(\U1761/y[1] ), .a(\U1761/x[3] ), .b(
        \U1761/x[2] ), .c(\U1761/x[3] ), .d(\U1761/U30/Z ), .e(\U1761/x[2] ), 
        .f(\U1761/U30/Z ) );
    inv_1 \U1761/U30/U30/Uinv  ( .x(\U1761/U30/Z ), .a(\U1761/y[1] ) );
    aoi222_1 \U1761/U31/U30/U1  ( .x(\U1761/x[1] ), .a(\nchdr_ack[3] ), .b(
        \nchdr_ack[2] ), .c(\nchdr_ack[3] ), .d(\U1761/U31/Z ), .e(
        \nchdr_ack[2] ), .f(\U1761/U31/Z ) );
    inv_1 \U1761/U31/U30/Uinv  ( .x(\U1761/U31/Z ), .a(\U1761/x[1] ) );
    aoi222_1 \U1632/U30/U1  ( .x(net178), .a(cack), .b(chdrctrlack), .c(cack), 
        .d(\U1632/Z ), .e(chdrctrlack), .f(\U1632/Z ) );
    inv_1 \U1632/U30/Uinv  ( .x(\U1632/Z ), .a(net178) );
    aoi222_1 \U1676/U30/U1  ( .x(hdrcd), .a(\chdrack[0] ), .b(\chdrack[1] ), 
        .c(\chdrack[0] ), .d(\U1676/Z ), .e(\chdrack[1] ), .f(\U1676/Z ) );
    inv_1 \U1676/U30/Uinv  ( .x(\U1676/Z ), .a(hdrcd) );
    nor3_1 \U1770/U21/Unr  ( .x(\U1770/U21/nr ), .a(\nchdr_ack[10] ), .b(
        \nchdr_ack[9] ), .c(\nchdr_ack[8] ) );
    nand3_1 \U1770/U21/Und  ( .x(\U1770/U21/nd ), .a(\nchdr_ack[10] ), .b(
        \nchdr_ack[9] ), .c(\nchdr_ack[8] ) );
    oa21_1 \U1770/U21/U1  ( .x(\U1770/U21/n2 ), .a(\U1770/U21/n2 ), .b(
        \U1770/U21/nr ), .c(\U1770/U21/nd ) );
    inv_1 \U1770/U21/U3  ( .x(\chdrack[1] ), .a(\U1770/U21/n2 ) );
    nor2_1 \U1652_0_/U2/U5  ( .x(\nchdr_ack[0] ), .a(\net242[10] ), .b(
        \net244[10] ) );
    ao222_2 \U1652_0_/U12/U19/U1/U1  ( .x(\net244[10] ), .a(\net243[10] ), .b(
        csize[0]), .c(\net243[10] ), .d(\net244[10] ), .e(csize[0]), .f(
        \net244[10] ) );
    ao222_2 \U1652_0_/U11/U19/U1/U1  ( .x(\net242[10] ), .a(csize[2]), .b(
        \net243[10] ), .c(csize[2]), .d(\net242[10] ), .e(\net243[10] ), .f(
        \net242[10] ) );
    nor2_1 \U1652_1_/U2/U5  ( .x(\nchdr_ack[1] ), .a(\net242[9] ), .b(
        \net244[9] ) );
    ao222_2 \U1652_1_/U12/U19/U1/U1  ( .x(\net244[9] ), .a(\net243[9] ), .b(
        csize[1]), .c(\net243[9] ), .d(\net244[9] ), .e(csize[1]), .f(
        \net244[9] ) );
    ao222_2 \U1652_1_/U11/U19/U1/U1  ( .x(\net242[9] ), .a(csize[3]), .b(
        \net243[9] ), .c(csize[3]), .d(\net242[9] ), .e(\net243[9] ), .f(
        \net242[9] ) );
    nor2_1 \U1652_2_/U2/U5  ( .x(\nchdr_ack[2] ), .a(\net242[8] ), .b(
        \net244[8] ) );
    ao222_2 \U1652_2_/U12/U19/U1/U1  ( .x(\net244[8] ), .a(\net243[8] ), .b(
        crnw[0]), .c(\net243[8] ), .d(\net244[8] ), .e(crnw[0]), .f(
        \net244[8] ) );
    ao222_2 \U1652_2_/U11/U19/U1/U1  ( .x(\net242[8] ), .a(crnw[1]), .b(
        \net243[8] ), .c(crnw[1]), .d(\net242[8] ), .e(\net243[8] ), .f(
        \net242[8] ) );
    nor2_1 \U1652_3_/U2/U5  ( .x(\nchdr_ack[3] ), .a(\net242[7] ), .b(
        \net244[7] ) );
    ao222_2 \U1652_3_/U12/U19/U1/U1  ( .x(\net244[7] ), .a(\net243[7] ), .b(
        ctag[0]), .c(\net243[7] ), .d(\net244[7] ), .e(ctag[0]), .f(
        \net244[7] ) );
    ao222_2 \U1652_3_/U11/U19/U1/U1  ( .x(\net242[7] ), .a(ctag[5]), .b(
        \net243[7] ), .c(ctag[5]), .d(\net242[7] ), .e(\net243[7] ), .f(
        \net242[7] ) );
    nor2_1 \U1652_4_/U2/U5  ( .x(\nchdr_ack[4] ), .a(\net242[6] ), .b(
        \net244[6] ) );
    ao222_2 \U1652_4_/U12/U19/U1/U1  ( .x(\net244[6] ), .a(\net243[6] ), .b(
        ctag[1]), .c(\net243[6] ), .d(\net244[6] ), .e(ctag[1]), .f(
        \net244[6] ) );
    ao222_2 \U1652_4_/U11/U19/U1/U1  ( .x(\net242[6] ), .a(ctag[6]), .b(
        \net243[6] ), .c(ctag[6]), .d(\net242[6] ), .e(\net243[6] ), .f(
        \net242[6] ) );
    nor2_1 \U1652_5_/U2/U5  ( .x(\nchdr_ack[5] ), .a(\net242[5] ), .b(
        \net244[5] ) );
    ao222_2 \U1652_5_/U12/U19/U1/U1  ( .x(\net244[5] ), .a(\net243[5] ), .b(
        ctag[2]), .c(\net243[5] ), .d(\net244[5] ), .e(ctag[2]), .f(
        \net244[5] ) );
    ao222_2 \U1652_5_/U11/U19/U1/U1  ( .x(\net242[5] ), .a(ctag[7]), .b(
        \net243[5] ), .c(ctag[7]), .d(\net242[5] ), .e(\net243[5] ), .f(
        \net242[5] ) );
    nor2_1 \U1652_6_/U2/U5  ( .x(\nchdr_ack[6] ), .a(\net242[4] ), .b(
        \net244[4] ) );
    ao222_2 \U1652_6_/U12/U19/U1/U1  ( .x(\net244[4] ), .a(\net243[4] ), .b(
        ctag[3]), .c(\net243[4] ), .d(\net244[4] ), .e(ctag[3]), .f(
        \net244[4] ) );
    ao222_2 \U1652_6_/U11/U19/U1/U1  ( .x(\net242[4] ), .a(ctag[8]), .b(
        \net243[4] ), .c(ctag[8]), .d(\net242[4] ), .e(\net243[4] ), .f(
        \net242[4] ) );
    nor2_1 \U1652_7_/U2/U5  ( .x(\nchdr_ack[7] ), .a(\net242[3] ), .b(
        \net244[3] ) );
    ao222_2 \U1652_7_/U12/U19/U1/U1  ( .x(\net244[3] ), .a(\net243[3] ), .b(
        ctag[4]), .c(\net243[3] ), .d(\net244[3] ), .e(ctag[4]), .f(
        \net244[3] ) );
    ao222_2 \U1652_7_/U11/U19/U1/U1  ( .x(\net242[3] ), .a(ctag[9]), .b(
        \net243[3] ), .c(ctag[9]), .d(\net242[3] ), .e(\net243[3] ), .f(
        \net242[3] ) );
    nor2_1 \U1652_8_/U2/U5  ( .x(\nchdr_ack[8] ), .a(\net242[2] ), .b(
        \net244[2] ) );
    ao222_2 \U1652_8_/U12/U19/U1/U1  ( .x(\net244[2] ), .a(\net243[2] ), .b(
        ccol[0]), .c(\net243[2] ), .d(\net244[2] ), .e(ccol[0]), .f(
        \net244[2] ) );
    ao222_2 \U1652_8_/U11/U19/U1/U1  ( .x(\net242[2] ), .a(ccol[3]), .b(
        \net243[2] ), .c(ccol[3]), .d(\net242[2] ), .e(\net243[2] ), .f(
        \net242[2] ) );
    nor2_1 \U1652_9_/U2/U5  ( .x(\nchdr_ack[9] ), .a(\net242[1] ), .b(
        \net244[1] ) );
    ao222_2 \U1652_9_/U12/U19/U1/U1  ( .x(\net244[1] ), .a(\net243[1] ), .b(
        ccol[1]), .c(\net243[1] ), .d(\net244[1] ), .e(ccol[1]), .f(
        \net244[1] ) );
    ao222_2 \U1652_9_/U11/U19/U1/U1  ( .x(\net242[1] ), .a(ccol[4]), .b(
        \net243[1] ), .c(ccol[4]), .d(\net242[1] ), .e(\net243[1] ), .f(
        \net242[1] ) );
    nor2_1 \U1652_10_/U2/U5  ( .x(\nchdr_ack[10] ), .a(\net242[0] ), .b(
        \net244[0] ) );
    ao222_2 \U1652_10_/U12/U19/U1/U1  ( .x(\net244[0] ), .a(\net243[0] ), .b(
        ccol[2]), .c(\net243[0] ), .d(\net244[0] ), .e(ccol[2]), .f(
        \net244[0] ) );
    ao222_2 \U1652_10_/U11/U19/U1/U1  ( .x(\net242[0] ), .a(ccol[5]), .b(
        \net243[0] ), .c(ccol[5]), .d(\net242[0] ), .e(\net243[0] ), .f(
        \net242[0] ) );
    nor2_1 \U1574_0_/U2/U5  ( .x(\U1574_0_/net231 ), .a(\rhdr_l[5] ), .b(
        \rhdr_h[5] ) );
    and2_1 \U1574_0_/U13/U8  ( .x(\net243[10] ), .a(\U1574_0_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_0_/U12/U19/U1/U1  ( .x(\rhdr_h[5] ), .a(n10), .b(
        \net242[10] ), .c(n10), .d(\rhdr_h[5] ), .e(\net242[10] ), .f(
        \rhdr_h[5] ) );
    ao222_2 \U1574_0_/U11/U19/U1/U1  ( .x(\rhdr_l[5] ), .a(\net244[10] ), .b(
        n9), .c(\net244[10] ), .d(\rhdr_l[5] ), .e(n10), .f(\rhdr_l[5] ) );
    nor2_1 \U1574_1_/U2/U5  ( .x(\U1574_1_/net231 ), .a(\rhdr_l[6] ), .b(
        \rhdr_h[6] ) );
    and2_1 \U1574_1_/U13/U8  ( .x(\net243[9] ), .a(\U1574_1_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_1_/U12/U19/U1/U1  ( .x(\rhdr_h[6] ), .a(n9), .b(\net242[9] 
        ), .c(n8), .d(\rhdr_h[6] ), .e(\net242[9] ), .f(\rhdr_h[6] ) );
    ao222_2 \U1574_1_/U11/U19/U1/U1  ( .x(\rhdr_l[6] ), .a(\net244[9] ), .b(n9
        ), .c(\net244[9] ), .d(\rhdr_l[6] ), .e(n10), .f(\rhdr_l[6] ) );
    nor2_1 \U1574_2_/U2/U5  ( .x(\U1574_2_/net231 ), .a(\rhdr_l[7] ), .b(
        \rhdr_h[7] ) );
    and2_1 \U1574_2_/U13/U8  ( .x(\net243[8] ), .a(\U1574_2_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_2_/U12/U19/U1/U1  ( .x(\rhdr_h[7] ), .a(n8), .b(\net242[8] 
        ), .c(n8), .d(\rhdr_h[7] ), .e(\net242[8] ), .f(\rhdr_h[7] ) );
    ao222_2 \U1574_2_/U11/U19/U1/U1  ( .x(\rhdr_l[7] ), .a(\net244[8] ), .b(n9
        ), .c(\net244[8] ), .d(\rhdr_l[7] ), .e(n10), .f(\rhdr_l[7] ) );
    nor2_1 \U1574_3_/U2/U5  ( .x(\U1574_3_/net231 ), .a(tag_l[0]), .b(tag_h[0]
        ) );
    and2_1 \U1574_3_/U13/U8  ( .x(\net243[7] ), .a(\U1574_3_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_3_/U12/U19/U1/U1  ( .x(tag_h[0]), .a(n10), .b(\net242[7] ), 
        .c(n8), .d(tag_h[0]), .e(\net242[7] ), .f(tag_h[0]) );
    ao222_2 \U1574_3_/U11/U19/U1/U1  ( .x(tag_l[0]), .a(\net244[7] ), .b(n9), 
        .c(\net244[7] ), .d(tag_l[0]), .e(n8), .f(tag_l[0]) );
    nor2_1 \U1574_4_/U2/U5  ( .x(\U1574_4_/net231 ), .a(tag_l[1]), .b(tag_h[1]
        ) );
    and2_1 \U1574_4_/U13/U8  ( .x(\net243[6] ), .a(\U1574_4_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_4_/U12/U19/U1/U1  ( .x(tag_h[1]), .a(n8), .b(\net242[6] ), 
        .c(n8), .d(tag_h[1]), .e(\net242[6] ), .f(tag_h[1]) );
    ao222_2 \U1574_4_/U11/U19/U1/U1  ( .x(tag_l[1]), .a(\net244[6] ), .b(n9), 
        .c(\net244[6] ), .d(tag_l[1]), .e(n8), .f(tag_l[1]) );
    nor2_1 \U1574_5_/U2/U5  ( .x(\U1574_5_/net231 ), .a(tag_l[2]), .b(tag_h[2]
        ) );
    and2_1 \U1574_5_/U13/U8  ( .x(\net243[5] ), .a(\U1574_5_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_5_/U12/U19/U1/U1  ( .x(tag_h[2]), .a(n9), .b(\net242[5] ), 
        .c(n8), .d(tag_h[2]), .e(\net242[5] ), .f(tag_h[2]) );
    ao222_2 \U1574_5_/U11/U19/U1/U1  ( .x(tag_l[2]), .a(\net244[5] ), .b(n9), 
        .c(\net244[5] ), .d(tag_l[2]), .e(n10), .f(tag_l[2]) );
    nor2_1 \U1574_6_/U2/U5  ( .x(\U1574_6_/net231 ), .a(tag_l[3]), .b(tag_h[3]
        ) );
    and2_1 \U1574_6_/U13/U8  ( .x(\net243[4] ), .a(\U1574_6_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_6_/U12/U19/U1/U1  ( .x(tag_h[3]), .a(n8), .b(\net242[4] ), 
        .c(n10), .d(tag_h[3]), .e(\net242[4] ), .f(tag_h[3]) );
    ao222_2 \U1574_6_/U11/U19/U1/U1  ( .x(tag_l[3]), .a(\net244[4] ), .b(n9), 
        .c(\net244[4] ), .d(tag_l[3]), .e(n8), .f(tag_l[3]) );
    nor2_1 \U1574_7_/U2/U5  ( .x(\U1574_7_/net231 ), .a(tag_l[4]), .b(tag_h[4]
        ) );
    and2_1 \U1574_7_/U13/U8  ( .x(\net243[3] ), .a(\U1574_7_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_7_/U12/U19/U1/U1  ( .x(tag_h[4]), .a(n8), .b(\net242[3] ), 
        .c(n10), .d(tag_h[4]), .e(\net242[3] ), .f(tag_h[4]) );
    ao222_2 \U1574_7_/U11/U19/U1/U1  ( .x(tag_l[4]), .a(\net244[3] ), .b(n9), 
        .c(\net244[3] ), .d(tag_l[4]), .e(n8), .f(tag_l[4]) );
    nor2_1 \U1574_8_/U2/U5  ( .x(\U1574_8_/net231 ), .a(\rhdr_l[13] ), .b(
        \rhdr_h[13] ) );
    and2_1 \U1574_8_/U13/U8  ( .x(\net243[2] ), .a(\U1574_8_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_8_/U12/U19/U1/U1  ( .x(\rhdr_h[13] ), .a(n9), .b(
        \net242[2] ), .c(n10), .d(\rhdr_h[13] ), .e(\net242[2] ), .f(
        \rhdr_h[13] ) );
    ao222_2 \U1574_8_/U11/U19/U1/U1  ( .x(\rhdr_l[13] ), .a(\net244[2] ), .b(
        n9), .c(\net244[2] ), .d(\rhdr_l[13] ), .e(n8), .f(\rhdr_l[13] ) );
    nor2_1 \U1574_9_/U2/U5  ( .x(\U1574_9_/net231 ), .a(\rhdr_l[14] ), .b(
        \rhdr_h[14] ) );
    and2_1 \U1574_9_/U13/U8  ( .x(\net243[1] ), .a(\U1574_9_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_9_/U12/U19/U1/U1  ( .x(\rhdr_h[14] ), .a(n10), .b(
        \net242[1] ), .c(n8), .d(\rhdr_h[14] ), .e(\net242[1] ), .f(
        \rhdr_h[14] ) );
    ao222_2 \U1574_9_/U11/U19/U1/U1  ( .x(\rhdr_l[14] ), .a(\net244[1] ), .b(
        n9), .c(\net244[1] ), .d(\rhdr_l[14] ), .e(n10), .f(\rhdr_l[14] ) );
    nor2_1 \U1574_10_/U2/U5  ( .x(\U1574_10_/net231 ), .a(\rhdr_l[15] ), .b(
        \rhdr_h[15] ) );
    and2_1 \U1574_10_/U13/U8  ( .x(\net243[0] ), .a(\U1574_10_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_10_/U12/U19/U1/U1  ( .x(\rhdr_h[15] ), .a(n10), .b(
        \net242[0] ), .c(n10), .d(\rhdr_h[15] ), .e(\net242[0] ), .f(
        \rhdr_h[15] ) );
    ao222_2 \U1574_10_/U11/U19/U1/U1  ( .x(\rhdr_l[15] ), .a(\net244[0] ), .b(
        n9), .c(\net244[0] ), .d(\rhdr_l[15] ), .e(n10), .f(\rhdr_l[15] ) );
    buf_1 U1 ( .x(csize[0]), .a(n15) );
    buf_1 U2 ( .x(csize[1]), .a(n14) );
    buf_1 U3 ( .x(csize[3]), .a(n13) );
    inv_0 U4 ( .x(n4), .a(n12) );
    inv_2 U5 ( .x(crnw[0]), .a(n4) );
    buf_1 U6 ( .x(crnw[1]), .a(n11) );
    inv_5 U7 ( .x(n7), .a(net265) );
    buf_3 U8 ( .x(nbreset), .a(nReset) );
    buf_3 U9 ( .x(n8), .a(net248) );
    buf_3 U10 ( .x(n10), .a(net248) );
    buf_3 U11 ( .x(n9), .a(net248) );
    nor2_1 U12 ( .x(net248), .a(net265), .b(rhdrack) );
endmodule


module chain_selement_ga_1 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_12 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[1] , \c[0] ;
    chain_selement_ga_1 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_2 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_13 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[1] , \c[0] ;
    chain_selement_ga_2 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_3 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_14 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[1] , \c[0] , n1, n2;
    chain_selement_ga_3 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        n2), .e(n2) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(n2), .b(r[0]), .c(n2), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(n2), .b(r[1]), .c(n2), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
    inv_0 U1 ( .x(n1), .a(e[0]) );
    inv_2 U2 ( .x(n2), .a(n1) );
endmodule


module chain_selement_ga_74 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module resp_route_tx_wb ( o, rtxack, e_h, e_l, noa, r_h, r_l, rtxreq );
output [4:0] o;
input  [2:0] e_h;
input  [2:0] e_l;
input  [2:0] r_h;
input  [2:0] r_l;
input  noa, rtxreq;
output rtxack;
    wire \r2[2] , \r2[1] , \r2[0] , \r1[2] , \r1[1] , \r1[0] , \r0[2] , 
        \r0[1] , \r0[0] , \last[0] , \last[1] , \last[2] , \last[3] , 
        \net72[0] , \net72[1] , net56, net106, net103, eopsym, net87, net66, 
        net84, net77, \I8/nb , \I8/na , \I11/n5 , \I11/n1 , \I11/n2 , \I11/n3 , 
        \I11/n4 , \I7_0_/U25/U1/clr , \I7_0_/U25/U1/ob , \I7_1_/U25/U1/clr , 
        \I7_1_/U25/U1/ob ;
    assign o[3] = 1'b0;
    assign o[2] = 1'b0;
    chain_selement_ga_74 I9 ( .Aa(\last[0] ), .Br(eopsym), .Ar(net87), .Ba(
        net66) );
    route_symbol_13 I2 ( .o({\r1[2] , \r1[1] , \r1[0] }), .txack(net84), 
        .txack_last(\last[2] ), .e({e_h[1], e_l[1]}), .oa(net66), .r({r_h[1], 
        r_l[1]}), .txreq(net77) );
    route_symbol_14 I3 ( .o({\r0[2] , \r0[1] , \r0[0] }), .txack(net87), 
        .txack_last(\last[1] ), .e({e_h[0], e_l[0]}), .oa(net66), .r({r_h[0], 
        r_l[0]}), .txreq(net84) );
    route_symbol_12 I1 ( .o({\r2[2] , \r2[1] , \r2[0] }), .txack(net77), 
        .txack_last(\last[3] ), .e({e_h[2], e_l[2]}), .oa(net66), .r({r_h[2], 
        r_l[2]}), .txreq(rtxreq) );
    nor2_1 \I5/U5  ( .x(net106), .a(eopsym), .b(\r2[2] ) );
    nor2_1 \I16/U5  ( .x(net103), .a(\r1[2] ), .b(\r0[2] ) );
    or2_1 \I14_0_/U12  ( .x(\net72[1] ), .a(\r2[0] ), .b(\r1[0] ) );
    or2_1 \I14_1_/U12  ( .x(\net72[0] ), .a(\r2[1] ), .b(\r1[1] ) );
    nor3_1 \I8/U27  ( .x(\I8/nb ), .a(o[4]), .b(o[3]), .c(o[2]) );
    nor2_1 \I8/U26  ( .x(\I8/na ), .a(o[1]), .b(o[0]) );
    nand2_2 \I8/U29  ( .x(net66), .a(\I8/nb ), .b(\I8/na ) );
    and4_1 \I11/U16  ( .x(\I11/n5 ), .a(\I11/n1 ), .b(\I11/n2 ), .c(\I11/n3 ), 
        .d(\I11/n4 ) );
    inv_1 \I11/U1  ( .x(\I11/n1 ), .a(\last[3] ) );
    inv_1 \I11/U2  ( .x(\I11/n2 ), .a(\last[2] ) );
    inv_1 \I11/U3  ( .x(\I11/n3 ), .a(\last[1] ) );
    inv_1 \I11/U4  ( .x(\I11/n4 ), .a(\last[0] ) );
    inv_1 \I11/U5  ( .x(rtxack), .a(\I11/n5 ) );
    nand2_1 \I17/U5  ( .x(net56), .a(net106), .b(net103) );
    ao222_1 \I15/U18/U1/U1  ( .x(o[4]), .a(noa), .b(net56), .c(noa), .d(o[4]), 
        .e(net56), .f(o[4]) );
    oa31_1 \I7_0_/U25/U1/Uclr  ( .x(\I7_0_/U25/U1/clr ), .a(noa), .b(\r0[0] ), 
        .c(\net72[1] ), .d(o[0]) );
    oaoi211_1 \I7_0_/U25/U1/Uaoi  ( .x(\I7_0_/U25/U1/ob ), .a(\r0[0] ), .b(
        \net72[1] ), .c(noa), .d(\I7_0_/U25/U1/clr ) );
    inv_2 \I7_0_/U25/U1/Ui  ( .x(o[0]), .a(\I7_0_/U25/U1/ob ) );
    oa31_1 \I7_1_/U25/U1/Uclr  ( .x(\I7_1_/U25/U1/clr ), .a(noa), .b(\r0[1] ), 
        .c(\net72[0] ), .d(o[1]) );
    oaoi211_1 \I7_1_/U25/U1/Uaoi  ( .x(\I7_1_/U25/U1/ob ), .a(\r0[1] ), .b(
        \net72[0] ), .c(noa), .d(\I7_1_/U25/U1/clr ) );
    inv_2 \I7_1_/U25/U1/Ui  ( .x(o[1]), .a(\I7_1_/U25/U1/ob ) );
endmodule


module matched_delay_cp2slave_resp_wb ( x, a );
input  a;
output x;
    buf_1 I1 ( .x(x), .a(a) );
endmodule


module matched_delay_cp2slave_com_wb ( x, a );
input  a;
output x;
    buf_1 I1 ( .x(x), .a(a) );
endmodule


module sr2dr_word_6 ( i, req, h, l );
input  [31:0] i;
output [31:0] h;
output [31:0] l;
input  req;
    wire \U31/nl , \U31/ni , \U31/nh , \U30/nl , \U30/ni , \U30/nh , \U29/nl , 
        \U29/ni , \U29/nh , \U28/nl , \U28/ni , \U28/nh , \U27/nl , \U27/ni , 
        \U27/nh , \U26/nl , \U26/ni , \U26/nh , \U25/nl , \U25/ni , \U25/nh , 
        \U24/nl , \U24/ni , \U24/nh , \U23/nl , \U23/ni , \U23/nh , \U22/nl , 
        \U22/ni , \U22/nh , \U21/nl , \U21/ni , \U21/nh , \U20/nl , \U20/ni , 
        \U20/nh , \U19/nl , \U19/ni , \U19/nh , \U18/nl , \U18/ni , \U18/nh , 
        \U17/nl , \U17/ni , \U17/nh , \U16/nl , \U16/ni , \U16/nh , \U15/nl , 
        \U15/ni , \U15/nh , \U14/nl , \U14/ni , \U14/nh , \U13/nl , \U13/ni , 
        \U13/nh , \U12/nl , \U12/ni , \U12/nh , \U11/nl , \U11/ni , \U11/nh , 
        \U10/nl , \U10/ni , \U10/nh , \U9/nl , \U9/ni , \U9/nh , \U8/nl , 
        \U8/ni , \U8/nh , \U7/nl , \U7/ni , \U7/nh , \U6/nl , \U6/ni , \U6/nh , 
        \U5/nl , \U5/ni , \U5/nh , \U4/nl , \U4/ni , \U4/nh , \U3/nl , \U3/ni , 
        \U3/nh , \U2/nl , \U2/ni , \U2/nh , \U1/nl , \U1/ni , \U1/nh , \U0/nl , 
        \U0/ni , \U0/nh , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
    inv_1 \U31/Uii  ( .x(\U31/ni ), .a(i[31]) );
    inv_1 \U31/Uih  ( .x(\U31/nh ), .a(h[31]) );
    inv_1 \U31/Uil  ( .x(\U31/nl ), .a(l[31]) );
    ao23_1 \U31/Ucl/U1/U1  ( .x(l[31]), .a(n9), .b(l[31]), .c(n1), .d(\U31/ni 
        ), .e(\U31/nh ) );
    ao23_1 \U31/Uch/U1/U1  ( .x(h[31]), .a(n9), .b(h[31]), .c(n2), .d(i[31]), 
        .e(\U31/nl ) );
    inv_1 \U30/Uii  ( .x(\U30/ni ), .a(i[30]) );
    inv_1 \U30/Uih  ( .x(\U30/nh ), .a(h[30]) );
    inv_1 \U30/Uil  ( .x(\U30/nl ), .a(l[30]) );
    ao23_1 \U30/Ucl/U1/U1  ( .x(l[30]), .a(n8), .b(l[30]), .c(n1), .d(\U30/ni 
        ), .e(\U30/nh ) );
    ao23_1 \U30/Uch/U1/U1  ( .x(h[30]), .a(n8), .b(h[30]), .c(n1), .d(i[30]), 
        .e(\U30/nl ) );
    inv_1 \U29/Uii  ( .x(\U29/ni ), .a(i[29]) );
    inv_1 \U29/Uih  ( .x(\U29/nh ), .a(h[29]) );
    inv_1 \U29/Uil  ( .x(\U29/nl ), .a(l[29]) );
    ao23_1 \U29/Ucl/U1/U1  ( .x(l[29]), .a(n8), .b(l[29]), .c(n1), .d(\U29/ni 
        ), .e(\U29/nh ) );
    ao23_1 \U29/Uch/U1/U1  ( .x(h[29]), .a(n8), .b(h[29]), .c(n2), .d(i[29]), 
        .e(\U29/nl ) );
    inv_1 \U28/Uii  ( .x(\U28/ni ), .a(i[28]) );
    inv_1 \U28/Uih  ( .x(\U28/nh ), .a(h[28]) );
    inv_1 \U28/Uil  ( .x(\U28/nl ), .a(l[28]) );
    ao23_1 \U28/Ucl/U1/U1  ( .x(l[28]), .a(n8), .b(l[28]), .c(n2), .d(\U28/ni 
        ), .e(\U28/nh ) );
    ao23_1 \U28/Uch/U1/U1  ( .x(h[28]), .a(n8), .b(h[28]), .c(n2), .d(i[28]), 
        .e(\U28/nl ) );
    inv_1 \U27/Uii  ( .x(\U27/ni ), .a(i[27]) );
    inv_1 \U27/Uih  ( .x(\U27/nh ), .a(h[27]) );
    inv_1 \U27/Uil  ( .x(\U27/nl ), .a(l[27]) );
    ao23_1 \U27/Ucl/U1/U1  ( .x(l[27]), .a(n8), .b(l[27]), .c(n2), .d(\U27/ni 
        ), .e(\U27/nh ) );
    ao23_1 \U27/Uch/U1/U1  ( .x(h[27]), .a(n8), .b(h[27]), .c(n2), .d(i[27]), 
        .e(\U27/nl ) );
    inv_1 \U26/Uii  ( .x(\U26/ni ), .a(i[26]) );
    inv_1 \U26/Uih  ( .x(\U26/nh ), .a(h[26]) );
    inv_1 \U26/Uil  ( .x(\U26/nl ), .a(l[26]) );
    ao23_1 \U26/Ucl/U1/U1  ( .x(l[26]), .a(n7), .b(l[26]), .c(n2), .d(\U26/ni 
        ), .e(\U26/nh ) );
    ao23_1 \U26/Uch/U1/U1  ( .x(h[26]), .a(n7), .b(h[26]), .c(n4), .d(i[26]), 
        .e(\U26/nl ) );
    inv_1 \U25/Uii  ( .x(\U25/ni ), .a(i[25]) );
    inv_1 \U25/Uih  ( .x(\U25/nh ), .a(h[25]) );
    inv_1 \U25/Uil  ( .x(\U25/nl ), .a(l[25]) );
    ao23_1 \U25/Ucl/U1/U1  ( .x(l[25]), .a(n7), .b(l[25]), .c(n4), .d(\U25/ni 
        ), .e(\U25/nh ) );
    ao23_1 \U25/Uch/U1/U1  ( .x(h[25]), .a(n7), .b(h[25]), .c(n4), .d(i[25]), 
        .e(\U25/nl ) );
    inv_1 \U24/Uii  ( .x(\U24/ni ), .a(i[24]) );
    inv_1 \U24/Uih  ( .x(\U24/nh ), .a(h[24]) );
    inv_1 \U24/Uil  ( .x(\U24/nl ), .a(l[24]) );
    ao23_1 \U24/Ucl/U1/U1  ( .x(l[24]), .a(n7), .b(l[24]), .c(n4), .d(\U24/ni 
        ), .e(\U24/nh ) );
    ao23_1 \U24/Uch/U1/U1  ( .x(h[24]), .a(n7), .b(h[24]), .c(n4), .d(i[24]), 
        .e(\U24/nl ) );
    inv_1 \U23/Uii  ( .x(\U23/ni ), .a(i[23]) );
    inv_1 \U23/Uih  ( .x(\U23/nh ), .a(h[23]) );
    inv_1 \U23/Uil  ( .x(\U23/nl ), .a(l[23]) );
    ao23_1 \U23/Ucl/U1/U1  ( .x(l[23]), .a(n7), .b(l[23]), .c(n3), .d(\U23/ni 
        ), .e(\U23/nh ) );
    ao23_1 \U23/Uch/U1/U1  ( .x(h[23]), .a(n7), .b(h[23]), .c(n3), .d(i[23]), 
        .e(\U23/nl ) );
    inv_1 \U22/Uii  ( .x(\U22/ni ), .a(i[22]) );
    inv_1 \U22/Uih  ( .x(\U22/nh ), .a(h[22]) );
    inv_1 \U22/Uil  ( .x(\U22/nl ), .a(l[22]) );
    ao23_1 \U22/Ucl/U1/U1  ( .x(l[22]), .a(n6), .b(l[22]), .c(n3), .d(\U22/ni 
        ), .e(\U22/nh ) );
    ao23_1 \U22/Uch/U1/U1  ( .x(h[22]), .a(n6), .b(h[22]), .c(n3), .d(i[22]), 
        .e(\U22/nl ) );
    inv_1 \U21/Uii  ( .x(\U21/ni ), .a(i[21]) );
    inv_1 \U21/Uih  ( .x(\U21/nh ), .a(h[21]) );
    inv_1 \U21/Uil  ( .x(\U21/nl ), .a(l[21]) );
    ao23_1 \U21/Ucl/U1/U1  ( .x(l[21]), .a(n6), .b(l[21]), .c(n3), .d(\U21/ni 
        ), .e(\U21/nh ) );
    ao23_1 \U21/Uch/U1/U1  ( .x(h[21]), .a(n6), .b(h[21]), .c(n3), .d(i[21]), 
        .e(\U21/nl ) );
    inv_1 \U20/Uii  ( .x(\U20/ni ), .a(i[20]) );
    inv_1 \U20/Uih  ( .x(\U20/nh ), .a(h[20]) );
    inv_1 \U20/Uil  ( .x(\U20/nl ), .a(l[20]) );
    ao23_1 \U20/Ucl/U1/U1  ( .x(l[20]), .a(n6), .b(l[20]), .c(n5), .d(\U20/ni 
        ), .e(\U20/nh ) );
    ao23_1 \U20/Uch/U1/U1  ( .x(h[20]), .a(n6), .b(h[20]), .c(n4), .d(i[20]), 
        .e(\U20/nl ) );
    inv_1 \U19/Uii  ( .x(\U19/ni ), .a(i[19]) );
    inv_1 \U19/Uih  ( .x(\U19/nh ), .a(h[19]) );
    inv_1 \U19/Uil  ( .x(\U19/nl ), .a(l[19]) );
    ao23_1 \U19/Ucl/U1/U1  ( .x(l[19]), .a(n6), .b(l[19]), .c(n4), .d(\U19/ni 
        ), .e(\U19/nh ) );
    ao23_1 \U19/Uch/U1/U1  ( .x(h[19]), .a(n6), .b(h[19]), .c(n4), .d(i[19]), 
        .e(\U19/nl ) );
    inv_1 \U18/Uii  ( .x(\U18/ni ), .a(i[18]) );
    inv_1 \U18/Uih  ( .x(\U18/nh ), .a(h[18]) );
    inv_1 \U18/Uil  ( .x(\U18/nl ), .a(l[18]) );
    ao23_1 \U18/Ucl/U1/U1  ( .x(l[18]), .a(n5), .b(l[18]), .c(n5), .d(\U18/ni 
        ), .e(\U18/nh ) );
    ao23_1 \U18/Uch/U1/U1  ( .x(h[18]), .a(n5), .b(h[18]), .c(n5), .d(i[18]), 
        .e(\U18/nl ) );
    inv_1 \U17/Uii  ( .x(\U17/ni ), .a(i[17]) );
    inv_1 \U17/Uih  ( .x(\U17/nh ), .a(h[17]) );
    inv_1 \U17/Uil  ( .x(\U17/nl ), .a(l[17]) );
    ao23_1 \U17/Ucl/U1/U1  ( .x(l[17]), .a(n6), .b(l[17]), .c(n5), .d(\U17/ni 
        ), .e(\U17/nh ) );
    ao23_1 \U17/Uch/U1/U1  ( .x(h[17]), .a(n7), .b(h[17]), .c(n4), .d(i[17]), 
        .e(\U17/nl ) );
    inv_1 \U16/Uii  ( .x(\U16/ni ), .a(i[16]) );
    inv_1 \U16/Uih  ( .x(\U16/nh ), .a(h[16]) );
    inv_1 \U16/Uil  ( .x(\U16/nl ), .a(l[16]) );
    ao23_1 \U16/Ucl/U1/U1  ( .x(l[16]), .a(n9), .b(l[16]), .c(n3), .d(\U16/ni 
        ), .e(\U16/nh ) );
    ao23_1 \U16/Uch/U1/U1  ( .x(h[16]), .a(n9), .b(h[16]), .c(n1), .d(i[16]), 
        .e(\U16/nl ) );
    inv_1 \U15/Uii  ( .x(\U15/ni ), .a(i[15]) );
    inv_1 \U15/Uih  ( .x(\U15/nh ), .a(h[15]) );
    inv_1 \U15/Uil  ( .x(\U15/nl ), .a(l[15]) );
    ao23_1 \U15/Ucl/U1/U1  ( .x(l[15]), .a(n8), .b(l[15]), .c(n1), .d(\U15/ni 
        ), .e(\U15/nh ) );
    ao23_1 \U15/Uch/U1/U1  ( .x(h[15]), .a(n7), .b(h[15]), .c(n1), .d(i[15]), 
        .e(\U15/nl ) );
    inv_1 \U14/Uii  ( .x(\U14/ni ), .a(i[14]) );
    inv_1 \U14/Uih  ( .x(\U14/nh ), .a(h[14]) );
    inv_1 \U14/Uil  ( .x(\U14/nl ), .a(l[14]) );
    ao23_1 \U14/Ucl/U1/U1  ( .x(l[14]), .a(n6), .b(l[14]), .c(n1), .d(\U14/ni 
        ), .e(\U14/nh ) );
    ao23_1 \U14/Uch/U1/U1  ( .x(h[14]), .a(n6), .b(h[14]), .c(n3), .d(i[14]), 
        .e(\U14/nl ) );
    inv_1 \U13/Uii  ( .x(\U13/ni ), .a(i[13]) );
    inv_1 \U13/Uih  ( .x(\U13/nh ), .a(h[13]) );
    inv_1 \U13/Uil  ( .x(\U13/nl ), .a(l[13]) );
    ao23_1 \U13/Ucl/U1/U1  ( .x(l[13]), .a(n6), .b(l[13]), .c(n4), .d(\U13/ni 
        ), .e(\U13/nh ) );
    ao23_1 \U13/Uch/U1/U1  ( .x(h[13]), .a(n6), .b(h[13]), .c(n4), .d(i[13]), 
        .e(\U13/nl ) );
    inv_1 \U12/Uii  ( .x(\U12/ni ), .a(i[12]) );
    inv_1 \U12/Uih  ( .x(\U12/nh ), .a(h[12]) );
    inv_1 \U12/Uil  ( .x(\U12/nl ), .a(l[12]) );
    ao23_1 \U12/Ucl/U1/U1  ( .x(l[12]), .a(n5), .b(l[12]), .c(n4), .d(\U12/ni 
        ), .e(\U12/nh ) );
    ao23_1 \U12/Uch/U1/U1  ( .x(h[12]), .a(n5), .b(h[12]), .c(n4), .d(i[12]), 
        .e(\U12/nl ) );
    inv_1 \U11/Uii  ( .x(\U11/ni ), .a(i[11]) );
    inv_1 \U11/Uih  ( .x(\U11/nh ), .a(h[11]) );
    inv_1 \U11/Uil  ( .x(\U11/nl ), .a(l[11]) );
    ao23_1 \U11/Ucl/U1/U1  ( .x(l[11]), .a(n5), .b(l[11]), .c(n4), .d(\U11/ni 
        ), .e(\U11/nh ) );
    ao23_1 \U11/Uch/U1/U1  ( .x(h[11]), .a(n5), .b(h[11]), .c(n4), .d(i[11]), 
        .e(\U11/nl ) );
    inv_1 \U10/Uii  ( .x(\U10/ni ), .a(i[10]) );
    inv_1 \U10/Uih  ( .x(\U10/nh ), .a(h[10]) );
    inv_1 \U10/Uil  ( .x(\U10/nl ), .a(l[10]) );
    ao23_1 \U10/Ucl/U1/U1  ( .x(l[10]), .a(n5), .b(l[10]), .c(n3), .d(\U10/ni 
        ), .e(\U10/nh ) );
    ao23_1 \U10/Uch/U1/U1  ( .x(h[10]), .a(n5), .b(h[10]), .c(n3), .d(i[10]), 
        .e(\U10/nl ) );
    inv_1 \U9/Uii  ( .x(\U9/ni ), .a(i[9]) );
    inv_1 \U9/Uih  ( .x(\U9/nh ), .a(h[9]) );
    inv_1 \U9/Uil  ( .x(\U9/nl ), .a(l[9]) );
    ao23_1 \U9/Ucl/U1/U1  ( .x(l[9]), .a(n5), .b(l[9]), .c(n3), .d(\U9/ni ), 
        .e(\U9/nh ) );
    ao23_1 \U9/Uch/U1/U1  ( .x(h[9]), .a(n5), .b(h[9]), .c(n3), .d(i[9]), .e(
        \U9/nl ) );
    inv_1 \U8/Uii  ( .x(\U8/ni ), .a(i[8]) );
    inv_1 \U8/Uih  ( .x(\U8/nh ), .a(h[8]) );
    inv_1 \U8/Uil  ( .x(\U8/nl ), .a(l[8]) );
    ao23_1 \U8/Ucl/U1/U1  ( .x(l[8]), .a(n5), .b(l[8]), .c(n3), .d(\U8/ni ), 
        .e(\U8/nh ) );
    ao23_1 \U8/Uch/U1/U1  ( .x(h[8]), .a(n5), .b(h[8]), .c(n3), .d(i[8]), .e(
        \U8/nl ) );
    inv_1 \U7/Uii  ( .x(\U7/ni ), .a(i[7]) );
    inv_1 \U7/Uih  ( .x(\U7/nh ), .a(h[7]) );
    inv_1 \U7/Uil  ( .x(\U7/nl ), .a(l[7]) );
    ao23_1 \U7/Ucl/U1/U1  ( .x(l[7]), .a(n7), .b(l[7]), .c(n3), .d(\U7/ni ), 
        .e(\U7/nh ) );
    ao23_1 \U7/Uch/U1/U1  ( .x(h[7]), .a(n7), .b(h[7]), .c(n2), .d(i[7]), .e(
        \U7/nl ) );
    inv_1 \U6/Uii  ( .x(\U6/ni ), .a(i[6]) );
    inv_1 \U6/Uih  ( .x(\U6/nh ), .a(h[6]) );
    inv_1 \U6/Uil  ( .x(\U6/nl ), .a(l[6]) );
    ao23_1 \U6/Ucl/U1/U1  ( .x(l[6]), .a(n7), .b(l[6]), .c(n2), .d(\U6/ni ), 
        .e(\U6/nh ) );
    ao23_1 \U6/Uch/U1/U1  ( .x(h[6]), .a(n7), .b(h[6]), .c(n2), .d(i[6]), .e(
        \U6/nl ) );
    inv_1 \U5/Uii  ( .x(\U5/ni ), .a(i[5]) );
    inv_1 \U5/Uih  ( .x(\U5/nh ), .a(h[5]) );
    inv_1 \U5/Uil  ( .x(\U5/nl ), .a(l[5]) );
    ao23_1 \U5/Ucl/U1/U1  ( .x(l[5]), .a(n7), .b(l[5]), .c(n2), .d(\U5/ni ), 
        .e(\U5/nh ) );
    ao23_1 \U5/Uch/U1/U1  ( .x(h[5]), .a(n7), .b(h[5]), .c(n2), .d(i[5]), .e(
        \U5/nl ) );
    inv_1 \U4/Uii  ( .x(\U4/ni ), .a(i[4]) );
    inv_1 \U4/Uih  ( .x(\U4/nh ), .a(h[4]) );
    inv_1 \U4/Uil  ( .x(\U4/nl ), .a(l[4]) );
    ao23_1 \U4/Ucl/U1/U1  ( .x(l[4]), .a(n6), .b(l[4]), .c(n2), .d(\U4/ni ), 
        .e(\U4/nh ) );
    ao23_1 \U4/Uch/U1/U1  ( .x(h[4]), .a(n6), .b(h[4]), .c(n2), .d(i[4]), .e(
        \U4/nl ) );
    inv_1 \U3/Uii  ( .x(\U3/ni ), .a(i[3]) );
    inv_1 \U3/Uih  ( .x(\U3/nh ), .a(h[3]) );
    inv_1 \U3/Uil  ( .x(\U3/nl ), .a(l[3]) );
    ao23_1 \U3/Ucl/U1/U1  ( .x(l[3]), .a(n6), .b(l[3]), .c(n2), .d(\U3/ni ), 
        .e(\U3/nh ) );
    ao23_1 \U3/Uch/U1/U1  ( .x(h[3]), .a(n8), .b(h[3]), .c(n1), .d(i[3]), .e(
        \U3/nl ) );
    inv_1 \U2/Uii  ( .x(\U2/ni ), .a(i[2]) );
    inv_1 \U2/Uih  ( .x(\U2/nh ), .a(h[2]) );
    inv_1 \U2/Uil  ( .x(\U2/nl ), .a(l[2]) );
    ao23_1 \U2/Ucl/U1/U1  ( .x(l[2]), .a(n8), .b(l[2]), .c(n1), .d(\U2/ni ), 
        .e(\U2/nh ) );
    ao23_1 \U2/Uch/U1/U1  ( .x(h[2]), .a(n8), .b(h[2]), .c(n1), .d(i[2]), .e(
        \U2/nl ) );
    inv_1 \U1/Uii  ( .x(\U1/ni ), .a(i[1]) );
    inv_1 \U1/Uih  ( .x(\U1/nh ), .a(h[1]) );
    inv_1 \U1/Uil  ( .x(\U1/nl ), .a(l[1]) );
    ao23_1 \U1/Ucl/U1/U1  ( .x(l[1]), .a(n8), .b(l[1]), .c(n1), .d(\U1/ni ), 
        .e(\U1/nh ) );
    ao23_1 \U1/Uch/U1/U1  ( .x(h[1]), .a(n8), .b(h[1]), .c(n1), .d(i[1]), .e(
        \U1/nl ) );
    inv_1 \U0/Uii  ( .x(\U0/ni ), .a(i[0]) );
    inv_1 \U0/Uih  ( .x(\U0/nh ), .a(h[0]) );
    inv_1 \U0/Uil  ( .x(\U0/nl ), .a(l[0]) );
    ao23_1 \U0/Ucl/U1/U1  ( .x(l[0]), .a(n8), .b(l[0]), .c(n1), .d(\U0/ni ), 
        .e(\U0/nh ) );
    ao23_1 \U0/Uch/U1/U1  ( .x(h[0]), .a(n8), .b(h[0]), .c(n1), .d(i[0]), .e(
        \U0/nl ) );
    buf_16 U1 ( .x(n1), .a(n12) );
    buf_16 U2 ( .x(n2), .a(n12) );
    buf_16 U3 ( .x(n3), .a(n12) );
    buf_16 U4 ( .x(n4), .a(n11) );
    buf_16 U5 ( .x(n5), .a(n11) );
    buf_16 U6 ( .x(n6), .a(n11) );
    buf_16 U7 ( .x(n7), .a(n10) );
    buf_16 U8 ( .x(n8), .a(n10) );
    buf_16 U9 ( .x(n9), .a(n10) );
    buf_16 U10 ( .x(n10), .a(req) );
    buf_16 U11 ( .x(n11), .a(req) );
    buf_16 U12 ( .x(n12), .a(req) );
endmodule


module cp2slave_wb ( tc_seq, tc_size, tc_itag, tc_wd, tc_lock, tc_a, tc_rnw, 
    tc_ok, tc_defer, tc_slow, tc_ack, req_in, ts_i, st_i, we_i, mult_i, adr_i, 
    dat_i, seq_i, prd_i, sel_i, ack_in, tr_rd, tr_err, tr_size, tr_ack, tr_rnw, 
    req_out, dat_o, err_o, rty_o, acc_o, sel_o, mult_o, rt_o, ack_out, reset
     );
input  [1:0] tc_seq;
input  [3:0] tc_size;
input  [9:0] tc_itag;
input  [63:0] tc_wd;
input  [1:0] tc_lock;
input  [63:0] tc_a;
input  [1:0] tc_rnw;
output [2:0] ts_i;
output [4:0] st_i;
output [31:0] adr_i;
output [31:0] dat_i;
output [3:0] sel_i;
output [63:0] tr_rd;
output [1:0] tr_err;
output [3:0] tr_size;
output [1:0] tr_rnw;
input  [31:0] dat_o;
input  [3:0] sel_o;
input  [4:0] rt_o;
input  ack_in, tr_ack, req_out, err_o, rty_o, acc_o, mult_o, reset;
output tc_ok, tc_defer, tc_slow, tc_ack, req_in, we_i, mult_i, seq_i, prd_i, 
    ack_out;
    wire \tc_a[60] , \tc_a[58] , \tc_wd[63] , \tc_wd[62] , \tc_wd[61] , 
        \tc_wd[60] , \tc_wd[59] , \tc_wd[58] , \tc_wd[56] , \tc_wd[55] , 
        \tc_wd[54] , \tc_wd[53] , \tc_wd[52] , \tc_wd[51] , \tc_wd[50] , 
        \tc_wd[49] , \tc_wd[48] , \tc_wd[47] , \tc_wd[46] , \tc_wd[45] , 
        \tc_wd[44] , \tc_wd[43] , \tc_wd[40] , \tc_wd[39] , \tc_wd[38] , 
        \tc_wd[36] , \tc_wd[32] , \sel_i[2] , n121, n122, n123, n124, n125, 
        n126, n127, n128, n129, n130, n135, n136, n137, n141, n142, n180, n181, 
        n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, 
        n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, 
        n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, 
        n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
        n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, 
        n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, 
        n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, 
        n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, 
        n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, 
        n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, 
        n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, 
        n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, 
        n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, 
        n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, 
        n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, 
        n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, 
        n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, 
        n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, 
        n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
        n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
        n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
        n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
        n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
        n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
        n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
        n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
        n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
        n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
        n518, n519, n520, n521, n522, n523, n524, n525, n529, n530, n531, n532, 
        n3, n4, n5, complb1, complb0, comp_basic, complw1, complw0, comp_wd, 
        all_w, all_r, respond, _24_net_, _25_net_, _26_net_, req_out_delayed, 
        req_in_i, \cg_all_w/__tmp99/loop , \Usze1/nl , \Usze1/ni , \Usze1/nh , 
        \Usze0/nl , \Usze0/ni , \Usze0/nh , \Urnw/nl , \Urnw/ni , \Urnw/nh , 
        \Uerr/nl , \Uerr/ni , \Uerr/nh , n1, n2;
    assign \tc_wd[63]  = tc_wd[63];
    assign \tc_wd[62]  = tc_wd[62];
    assign \tc_wd[61]  = tc_wd[61];
    assign \tc_wd[60]  = tc_wd[60];
    assign \tc_wd[59]  = tc_wd[59];
    assign \tc_wd[58]  = tc_wd[58];
    assign \tc_wd[56]  = tc_wd[56];
    assign \tc_wd[55]  = tc_wd[55];
    assign \tc_wd[54]  = tc_wd[54];
    assign \tc_wd[53]  = tc_wd[53];
    assign \tc_wd[52]  = tc_wd[52];
    assign \tc_wd[51]  = tc_wd[51];
    assign \tc_wd[50]  = tc_wd[50];
    assign \tc_wd[49]  = tc_wd[49];
    assign \tc_wd[48]  = tc_wd[48];
    assign \tc_wd[47]  = tc_wd[47];
    assign \tc_wd[46]  = tc_wd[46];
    assign \tc_wd[45]  = tc_wd[45];
    assign \tc_wd[44]  = tc_wd[44];
    assign \tc_wd[43]  = tc_wd[43];
    assign \tc_wd[40]  = tc_wd[40];
    assign \tc_wd[39]  = tc_wd[39];
    assign \tc_wd[38]  = tc_wd[38];
    assign \tc_wd[36]  = tc_wd[36];
    assign \tc_wd[32]  = tc_wd[32];
    assign \tc_a[60]  = tc_a[60];
    assign \tc_a[58]  = tc_a[58];
    assign ts_i[2] = 1'b0;
    assign ts_i[1] = 1'b0;
    assign ts_i[0] = 1'b0;
    assign adr_i[28] = \tc_a[60] ;
    assign adr_i[26] = \tc_a[58] ;
    assign dat_i[31] = \tc_wd[63] ;
    assign dat_i[30] = \tc_wd[62] ;
    assign dat_i[29] = \tc_wd[61] ;
    assign dat_i[28] = \tc_wd[60] ;
    assign dat_i[27] = \tc_wd[59] ;
    assign dat_i[26] = \tc_wd[58] ;
    assign dat_i[24] = \tc_wd[56] ;
    assign dat_i[23] = \tc_wd[55] ;
    assign dat_i[22] = \tc_wd[54] ;
    assign dat_i[21] = \tc_wd[53] ;
    assign dat_i[20] = \tc_wd[52] ;
    assign dat_i[19] = \tc_wd[51] ;
    assign dat_i[18] = \tc_wd[50] ;
    assign dat_i[17] = \tc_wd[49] ;
    assign dat_i[16] = \tc_wd[48] ;
    assign dat_i[15] = \tc_wd[47] ;
    assign dat_i[14] = \tc_wd[46] ;
    assign dat_i[13] = \tc_wd[45] ;
    assign dat_i[12] = \tc_wd[44] ;
    assign dat_i[11] = \tc_wd[43] ;
    assign dat_i[8] = \tc_wd[40] ;
    assign dat_i[7] = \tc_wd[39] ;
    assign dat_i[6] = \tc_wd[38] ;
    assign dat_i[4] = \tc_wd[36] ;
    assign dat_i[0] = \tc_wd[32] ;
    assign prd_i = 1'b0;
    assign sel_i[3] = \sel_i[2] ;
    assign sel_i[2] = \sel_i[2] ;
    assign sel_i[0] = 1'b1;
    assign tc_ack = ack_in;
    assign ack_out = tr_ack;
    sr2dr_word_6 Urd ( .i(dat_o), .req(n1), .h(tr_rd[63:32]), .l(tr_rd[31:0])
         );
    inv_1 U3 ( .x(n334), .a(tc_a[7]) );
    inv_1 U5 ( .x(n311), .a(tc_a[21]) );
    and2_1 U6 ( .x(n129), .a(n309), .b(n310) );
    inv_1 U7 ( .x(n309), .a(tc_a[6]) );
    inv_1 U9 ( .x(n315), .a(tc_itag[4]) );
    nand2_1 U10 ( .x(n348), .a(n349), .b(n350) );
    inv_1 U11 ( .x(n349), .a(tc_a[12]) );
    inv_1 U12 ( .x(n456), .a(n348) );
    inv_1 U13 ( .x(n336), .a(tc_a[30]) );
    inv_1 U14 ( .x(n457), .a(n345) );
    inv_1 U15 ( .x(n303), .a(tc_a[8]) );
    nand3_1 U16 ( .x(n505), .a(n193), .b(n476), .c(n479) );
    inv_1 U17 ( .x(n229), .a(tc_wd[5]) );
    inv_1 U18 ( .x(n226), .a(tc_wd[3]) );
    inv_1 U19 ( .x(n257), .a(tc_wd[16]) );
    inv_1 U20 ( .x(n263), .a(tc_wd[21]) );
    inv_1 U21 ( .x(n260), .a(tc_wd[19]) );
    nand2_1 U22 ( .x(n268), .a(n269), .b(n270) );
    inv_1 U23 ( .x(n269), .a(tc_wd[23]) );
    inv_1 U24 ( .x(n270), .a(\tc_wd[55] ) );
    nand2_1 U25 ( .x(n265), .a(n266), .b(n267) );
    inv_1 U26 ( .x(n266), .a(tc_wd[20]) );
    inv_1 U27 ( .x(n277), .a(tc_wd[27]) );
    inv_1 U28 ( .x(n252), .a(\tc_wd[47] ) );
    nand2_1 U29 ( .x(n248), .a(n249), .b(n250) );
    inv_1 U30 ( .x(n249), .a(tc_wd[12]) );
    nand2_1 U31 ( .x(n245), .a(n246), .b(n247) );
    inv_1 U32 ( .x(n246), .a(tc_wd[13]) );
    inv_1 U33 ( .x(n247), .a(\tc_wd[45] ) );
    nand2_1 U34 ( .x(n242), .a(n243), .b(n244) );
    inv_1 U35 ( .x(n243), .a(tc_wd[11]) );
    nand2_1 U36 ( .x(n222), .a(n223), .b(n224) );
    inv_1 U37 ( .x(n223), .a(tc_wd[0]) );
    inv_1 U38 ( .x(n220), .a(tc_wd[1]) );
    nand2_1 U39 ( .x(n234), .a(n235), .b(n236) );
    inv_1 U40 ( .x(n235), .a(tc_wd[7]) );
    nand2_1 U41 ( .x(n231), .a(n232), .b(n233) );
    inv_1 U42 ( .x(n232), .a(tc_wd[4]) );
    nand2_1 U43 ( .x(n205), .a(n206), .b(n207) );
    inv_1 U44 ( .x(n206), .a(tc_wd[18]) );
    inv_1 U45 ( .x(n203), .a(tc_wd[10]) );
    nand2_1 U46 ( .x(n199), .a(n200), .b(n201) );
    inv_1 U47 ( .x(n200), .a(tc_wd[6]) );
    inv_1 U48 ( .x(n197), .a(tc_wd[2]) );
    inv_1 U49 ( .x(n218), .a(\tc_wd[46] ) );
    nand2_1 U50 ( .x(n214), .a(n215), .b(n216) );
    inv_1 U51 ( .x(n215), .a(tc_wd[30]) );
    nand2_1 U52 ( .x(n211), .a(n212), .b(n213) );
    inv_1 U53 ( .x(n213), .a(\tc_wd[58] ) );
    nand2_1 U54 ( .x(n208), .a(n209), .b(n210) );
    inv_1 U55 ( .x(n209), .a(tc_wd[22]) );
    inv_1 U56 ( .x(n374), .a(tc_rnw[0]) );
    inv_1 U57 ( .x(n375), .a(tc_rnw[1]) );
    inv_1 U58 ( .x(n368), .a(tc_a[18]) );
    inv_1 U59 ( .x(n244), .a(\tc_wd[43] ) );
    inv_1 U60 ( .x(n251), .a(tc_wd[15]) );
    inv_1 U61 ( .x(n250), .a(\tc_wd[44] ) );
    inv_1 U62 ( .x(n280), .a(tc_wd[29]) );
    inv_1 U63 ( .x(n267), .a(\tc_wd[52] ) );
    inv_1 U64 ( .x(n274), .a(tc_wd[24]) );
    inv_1 U65 ( .x(n271), .a(tc_wd[25]) );
    inv_1 U66 ( .x(n212), .a(tc_wd[26]) );
    inv_1 U67 ( .x(n210), .a(\tc_wd[54] ) );
    inv_1 U68 ( .x(n216), .a(\tc_wd[62] ) );
    inv_1 U69 ( .x(n201), .a(\tc_wd[38] ) );
    inv_1 U70 ( .x(n427), .a(n196) );
    inv_1 U71 ( .x(n207), .a(\tc_wd[50] ) );
    inv_1 U72 ( .x(n424), .a(n202) );
    inv_1 U73 ( .x(n236), .a(\tc_wd[39] ) );
    inv_1 U74 ( .x(n233), .a(\tc_wd[36] ) );
    inv_1 U75 ( .x(n240), .a(tc_wd[8]) );
    inv_1 U76 ( .x(n237), .a(tc_wd[9]) );
    inv_1 U77 ( .x(n224), .a(\tc_wd[32] ) );
    inv_1 U78 ( .x(n413), .a(n219) );
    nand2_1 U79 ( .x(n421), .a(n418), .b(n416) );
    nand2_1 U80 ( .x(n428), .a(n425), .b(n422) );
    nand2_1 U81 ( .x(n414), .a(n411), .b(n408) );
    inv_1 U82 ( .x(n238), .a(tc_wd[41]) );
    inv_1 U83 ( .x(n272), .a(tc_wd[57]) );
    inv_1 U84 ( .x(n350), .a(tc_a[44]) );
    inv_1 U85 ( .x(n351), .a(tc_a[43]) );
    inv_1 U86 ( .x(n366), .a(tc_a[41]) );
    inv_1 U87 ( .x(n335), .a(tc_a[39]) );
    inv_1 U88 ( .x(n310), .a(tc_a[38]) );
    inv_1 U89 ( .x(n355), .a(tc_a[52]) );
    and3_1 U90 ( .x(tc_ok), .a(n531), .b(n532), .c(respond) );
    and2_1 U91 ( .x(tc_slow), .a(respond), .b(acc_o) );
    inv_1 U94 ( .x(n313), .a(tc_itag[5]) );
    and2_1 U95 ( .x(n121), .a(n334), .b(n335) );
    and2_1 U96 ( .x(n122), .a(n359), .b(n360) );
    and2_1 U97 ( .x(n123), .a(n336), .b(n337) );
    and2_1 U98 ( .x(n124), .a(n237), .b(n238) );
    and2_1 U99 ( .x(n125), .a(n251), .b(n252) );
    and2_1 U100 ( .x(n126), .a(n271), .b(n272) );
    and2_1 U101 ( .x(n127), .a(n217), .b(n218) );
    and2_1 U102 ( .x(n128), .a(n311), .b(n312) );
    nor2_1 U103 ( .x(n130), .a(tc_size[3]), .b(tc_size[2]) );
    nand2i_1 U105 ( .x(n284), .a(tc_wd[31]), .b(n285) );
    oa22_1 U106 ( .x(n449), .a(tc_a[27]), .b(tc_a[59]), .c(tc_a[54]), .d(tc_a
        [22]) );
    inv_1 U107 ( .x(n359), .a(tc_a[27]) );
    inv_1 U108 ( .x(n360), .a(tc_a[59]) );
    nand2i_1 U109 ( .x(n282), .a(tc_wd[28]), .b(n283) );
    nor2_1 U110 ( .x(n479), .a(tc_itag[0]), .b(tc_itag[5]) );
    nand4_1 U112 ( .x(n380), .a(n279), .b(n276), .c(n284), .d(n282) );
    aoi21_1 U113 ( .x(n425), .a(n200), .b(n201), .c(n427) );
    oa22_1 U114 ( .x(n397), .a(tc_wd[13]), .b(\tc_wd[45] ), .c(tc_wd[11]), .d(
        \tc_wd[43] ) );
    nor2_1 U115 ( .x(n454), .a(tc_a[20]), .b(tc_a[52]) );
    aoi21_1 U116 ( .x(n422), .a(n206), .b(n207), .c(n424) );
    oa22_1 U117 ( .x(n418), .a(tc_wd[26]), .b(\tc_wd[58] ), .c(tc_wd[22]), .d(
        \tc_wd[54] ) );
    oa22_1 U118 ( .x(n416), .a(tc_wd[14]), .b(\tc_wd[46] ), .c(tc_wd[30]), .d(
        \tc_wd[62] ) );
    inv_1 U119 ( .x(n217), .a(tc_wd[14]) );
    aoi22_1 U120 ( .x(n463), .a(n336), .b(n337), .c(n334), .d(n335) );
    nor2_1 U121 ( .x(n453), .a(tc_a[11]), .b(tc_a[43]) );
    oa22_1 U122 ( .x(n395), .a(tc_wd[15]), .b(\tc_wd[47] ), .c(tc_wd[12]), .d(
        \tc_wd[44] ) );
    oa22_1 U123 ( .x(n404), .a(tc_wd[7]), .b(\tc_wd[39] ), .c(tc_wd[4]), .d(
        \tc_wd[36] ) );
    oa22_1 U124 ( .x(n383), .a(tc_wd[23]), .b(\tc_wd[55] ), .c(tc_wd[20]), .d(
        \tc_wd[52] ) );
    aoi21_1 U125 ( .x(n411), .a(n223), .b(n224), .c(n413) );
    nor2_1 U126 ( .x(n443), .a(tc_a[49]), .b(tc_a[17]) );
    aoi22_1 U127 ( .x(n477), .a(n311), .b(n312), .c(n309), .d(n310) );
    oa21_1 U128 ( .x(n455), .a(tc_a[12]), .b(tc_a[44]), .c(n345) );
    inv_1 U129 ( .x(dat_i[5]), .a(n230) );
    inv_1 U130 ( .x(dat_i[9]), .a(n238) );
    inv_1 U131 ( .x(dat_i[25]), .a(n272) );
    buf_1 U132 ( .x(\sel_i[2] ), .a(tc_size[3]) );
    buf_1 U133 ( .x(adr_i[16]), .a(tc_a[48]) );
    nor2_1 U134 ( .x(n135), .a(tc_a[14]), .b(tc_a[46]) );
    inv_1 U135 ( .x(n305), .a(tc_a[46]) );
    inv_1 U136 ( .x(n487), .a(n302) );
    nand2i_1 U137 ( .x(n445), .a(n446), .b(n442) );
    nor2_1 U138 ( .x(n136), .a(tc_a[29]), .b(tc_a[61]) );
    inv_1 U139 ( .x(n320), .a(tc_a[61]) );
    nand2_1 U140 ( .x(n400), .a(n397), .b(n395) );
    inv_1 U141 ( .x(n137), .a(n340) );
    inv_1 U142 ( .x(dat_i[2]), .a(n198) );
    nand2_1 U143 ( .x(n386), .a(n383), .b(n381) );
    nand3i_1 U144 ( .x(n478), .a(n479), .b(n477), .c(n475) );
    nand2_1 U145 ( .x(n407), .a(n404), .b(n402) );
    inv_1 U146 ( .x(dat_i[10]), .a(n204) );
    inv_1 U147 ( .x(dat_i[1]), .a(n221) );
    nor2_1 U148 ( .x(n141), .a(tc_a[3]), .b(tc_a[35]) );
    inv_1 U149 ( .x(n321), .a(tc_a[35]) );
    nor2_1 U151 ( .x(n483), .a(n484), .b(n485) );
    nor2_1 U152 ( .x(n480), .a(n474), .b(n478) );
    inv_1 U153 ( .x(dat_i[3]), .a(n227) );
    nor2_1 U154 ( .x(n188), .a(n517), .b(n525) );
    nand2_1 U155 ( .x(n180), .a(n401), .b(n387) );
    nor2_1 U156 ( .x(n401), .a(n394), .b(n400) );
    nor2_1 U157 ( .x(n387), .a(n380), .b(n386) );
    nor2_1 U158 ( .x(n481), .a(n482), .b(n135) );
    nor2_1 U159 ( .x(n491), .a(n195), .b(n492) );
    nor2_1 U160 ( .x(n195), .a(tc_size[1]), .b(tc_size[3]) );
    inv_1 U161 ( .x(adr_i[18]), .a(n369) );
    nand2_1 U162 ( .x(n181), .a(n429), .b(n415) );
    nor2_1 U163 ( .x(n429), .a(n421), .b(n428) );
    nor2_1 U164 ( .x(n415), .a(n407), .b(n414) );
    inv_1 U165 ( .x(adr_i[0]), .a(n324) );
    inv_1 U166 ( .x(n324), .a(tc_a[32]) );
    inv_1 U167 ( .x(sel_i[1]), .a(n130) );
    inv_1 U168 ( .x(st_i[2]), .a(n343) );
    inv_1 U169 ( .x(adr_i[9]), .a(n366) );
    inv_1 U170 ( .x(adr_i[24]), .a(n363) );
    inv_1 U171 ( .x(adr_i[19]), .a(n319) );
    inv_1 U172 ( .x(n319), .a(tc_a[51]) );
    inv_1 U173 ( .x(n369), .a(tc_a[50]) );
    inv_1 U174 ( .x(st_i[3]), .a(n344) );
    inv_1 U175 ( .x(adr_i[13]), .a(n354) );
    inv_1 U176 ( .x(adr_i[12]), .a(n350) );
    inv_1 U177 ( .x(adr_i[8]), .a(n304) );
    inv_1 U178 ( .x(n304), .a(tc_a[40]) );
    inv_1 U179 ( .x(adr_i[2]), .a(n330) );
    buf_1 U180 ( .x(adr_i[17]), .a(tc_a[49]) );
    nand2_1 U181 ( .x(n497), .a(n496), .b(n130) );
    inv_1 U182 ( .x(adr_i[10]), .a(n291) );
    and2_1 U183 ( .x(n438), .a(n373), .b(n367) );
    inv_1 U184 ( .x(n439), .a(n373) );
    inv_1 U185 ( .x(n440), .a(n367) );
    inv_1 U186 ( .x(adr_i[20]), .a(n355) );
    inv_1 U187 ( .x(adr_i[27]), .a(n360) );
    inv_1 U188 ( .x(adr_i[4]), .a(n333) );
    inv_1 U189 ( .x(adr_i[25]), .a(n308) );
    inv_1 U190 ( .x(adr_i[30]), .a(n337) );
    inv_1 U191 ( .x(adr_i[31]), .a(n297) );
    inv_1 U192 ( .x(n297), .a(tc_a[63]) );
    inv_1 U193 ( .x(adr_i[15]), .a(n347) );
    inv_1 U194 ( .x(adr_i[11]), .a(n351) );
    inv_1 U195 ( .x(adr_i[1]), .a(n301) );
    inv_1 U196 ( .x(n301), .a(tc_a[33]) );
    nand2_1 U197 ( .x(n503), .a(n499), .b(n502) );
    nor2_1 U198 ( .x(n499), .a(n497), .b(n498) );
    inv_1 U199 ( .x(adr_i[21]), .a(n312) );
    inv_1 U200 ( .x(n312), .a(tc_a[53]) );
    inv_1 U201 ( .x(seq_i), .a(n288) );
    inv_1 U202 ( .x(adr_i[5]), .a(n327) );
    inv_1 U203 ( .x(st_i[4]), .a(n316) );
    inv_1 U204 ( .x(n316), .a(tc_itag[9]) );
    inv_1 U205 ( .x(st_i[1]), .a(n298) );
    inv_1 U206 ( .x(adr_i[23]), .a(n294) );
    inv_1 U207 ( .x(adr_i[22]), .a(n358) );
    nand2_1 U208 ( .x(complb0), .a(n188), .b(n189) );
    nor2_1 U209 ( .x(n189), .a(n503), .b(n510) );
    inv_1 U210 ( .x(adr_i[29]), .a(n320) );
    inv_1 U211 ( .x(adr_i[7]), .a(n335) );
    inv_1 U212 ( .x(adr_i[14]), .a(n305) );
    inv_1 U213 ( .x(adr_i[6]), .a(n310) );
    inv_1 U214 ( .x(st_i[0]), .a(n313) );
    inv_1 U215 ( .x(adr_i[3]), .a(n321) );
    nand3_1 U218 ( .x(n507), .a(n192), .b(n136), .c(n473) );
    nand2_1 U219 ( .x(n508), .a(n471), .b(n141) );
    nor2_1 U220 ( .x(n488), .a(n489), .b(n490) );
    nand4_1 U222 ( .x(complw0), .a(n182), .b(n183), .c(n184), .d(n185) );
    nor2_1 U223 ( .x(n192), .a(\tc_a[58] ), .b(tc_a[26]) );
    nor2_1 U224 ( .x(n193), .a(tc_a[48]), .b(tc_a[16]) );
    nand2_1 U225 ( .x(n364), .a(n365), .b(n366) );
    nand2_1 U226 ( .x(n394), .a(n391), .b(n388) );
    nand4_1 U227 ( .x(n430), .a(n423), .b(n424), .c(n426), .d(n427) );
    nand4_1 U228 ( .x(n431), .a(n127), .b(n417), .c(n419), .d(n420) );
    nor2_1 U229 ( .x(n185), .a(n430), .b(n431) );
    nand4_1 U230 ( .x(n432), .a(n409), .b(n410), .c(n412), .d(n413) );
    nand4_1 U231 ( .x(n433), .a(n403), .b(n124), .c(n405), .d(n406) );
    nor2_1 U232 ( .x(n184), .a(n432), .b(n433) );
    nand4_1 U233 ( .x(n434), .a(n125), .b(n396), .c(n398), .d(n399) );
    nand4_1 U234 ( .x(n435), .a(n389), .b(n390), .c(n392), .d(n393) );
    nor2_1 U235 ( .x(n183), .a(n434), .b(n435) );
    nand4_1 U236 ( .x(n436), .a(n382), .b(n126), .c(n384), .d(n385) );
    nand4_1 U237 ( .x(n437), .a(n376), .b(n377), .c(n378), .d(n379) );
    nor2_1 U238 ( .x(n182), .a(n436), .b(n437) );
    nand2_1 U239 ( .x(n441), .a(n438), .b(n370) );
    nor2_1 U240 ( .x(n442), .a(n443), .b(n444) );
    nor3_1 U241 ( .x(n470), .a(n471), .b(n136), .c(n141) );
    nor3_1 U242 ( .x(n472), .a(n473), .b(n192), .c(n193) );
    nand2_1 U243 ( .x(n474), .a(n472), .b(n470) );
    nor2_1 U244 ( .x(n475), .a(n476), .b(n194) );
    nand3i_1 U245 ( .x(n486), .a(n487), .b(n481), .c(n483) );
    nand3i_1 U246 ( .x(n493), .a(n494), .b(n488), .c(n491) );
    nor2_1 U247 ( .x(n495), .a(n493), .b(n486) );
    nand2_1 U248 ( .x(n191), .a(n495), .b(n480) );
    nand3_1 U249 ( .x(n498), .a(n489), .b(n492), .c(n490) );
    nand3_1 U250 ( .x(n500), .a(n485), .b(n494), .c(n484) );
    nand2_1 U251 ( .x(n501), .a(n135), .b(n487) );
    nor2_1 U252 ( .x(n502), .a(n500), .b(n501) );
    nand3_1 U253 ( .x(n504), .a(n128), .b(n482), .c(n129) );
    nor2_1 U254 ( .x(n506), .a(n504), .b(n505) );
    nor2_1 U255 ( .x(n509), .a(n507), .b(n508) );
    nand2_1 U256 ( .x(n510), .a(n509), .b(n506) );
    nand3_1 U257 ( .x(n511), .a(n465), .b(n466), .c(n468) );
    nand3_1 U258 ( .x(n512), .a(n123), .b(n121), .c(n460) );
    nor2_1 U259 ( .x(n513), .a(n511), .b(n512) );
    nand3_1 U260 ( .x(n514), .a(n462), .b(n459), .c(n457) );
    nand2_1 U261 ( .x(n515), .a(n453), .b(n456) );
    nor2_1 U262 ( .x(n516), .a(n514), .b(n515) );
    nand2_1 U263 ( .x(n517), .a(n516), .b(n513) );
    nand2_1 U264 ( .x(n518), .a(n454), .b(n452) );
    nor2i_1 U265 ( .x(n519), .a(n450), .b(n518) );
    nand2_1 U266 ( .x(n520), .a(n444), .b(n122) );
    nor2i_1 U267 ( .x(n522), .a(n446), .b(n521) );
    nand2_1 U268 ( .x(n523), .a(n439), .b(n524) );
    inv_1 U270 ( .x(n365), .a(tc_a[9]) );
    inv_1 U271 ( .x(n371), .a(\tc_a[60] ) );
    inv_1 U272 ( .x(n446), .a(n364) );
    nor2_1 U273 ( .x(complb1), .a(n190), .b(n191) );
    nor2_1 U274 ( .x(complw1), .a(n180), .b(n181) );
    nand3i_1 U276 ( .x(n190), .a(n441), .b(n447), .c(n469) );
    and4_1 U277 ( .x(n5), .a(n3), .b(n4), .c(n519), .d(n522) );
    inv_1 U216 ( .x(n3), .a(n520) );
    inv_1 U217 ( .x(n4), .a(n523) );
    inv_1 U428 ( .x(n525), .a(n5) );
    nor2_1 U278 ( .x(n447), .a(n448), .b(n445) );
    nor2_1 U279 ( .x(n469), .a(n467), .b(n461) );
    nand2_1 U280 ( .x(n370), .a(n371), .b(n372) );
    nand3i_1 U281 ( .x(n448), .a(n454), .b(n449), .c(n451) );
    nand3i_1 U282 ( .x(n461), .a(n462), .b(n455), .c(n458) );
    nand3i_1 U283 ( .x(n467), .a(n468), .b(n463), .c(n464) );
    inv_1 U284 ( .x(n382), .a(n273) );
    inv_1 U285 ( .x(n384), .a(n268) );
    inv_1 U286 ( .x(n385), .a(n265) );
    inv_1 U287 ( .x(n376), .a(n284) );
    inv_1 U288 ( .x(n377), .a(n282) );
    inv_1 U289 ( .x(n378), .a(n279) );
    inv_1 U290 ( .x(n379), .a(n276) );
    inv_1 U291 ( .x(n396), .a(n248) );
    inv_1 U292 ( .x(n398), .a(n245) );
    inv_1 U293 ( .x(n399), .a(n242) );
    inv_1 U294 ( .x(n389), .a(n262) );
    inv_1 U295 ( .x(n390), .a(n259) );
    inv_1 U296 ( .x(n392), .a(n256) );
    inv_1 U297 ( .x(n393), .a(n253) );
    inv_1 U298 ( .x(n409), .a(n228) );
    inv_1 U299 ( .x(n410), .a(n225) );
    inv_1 U300 ( .x(n412), .a(n222) );
    inv_1 U301 ( .x(n403), .a(n239) );
    inv_1 U302 ( .x(n405), .a(n234) );
    inv_1 U303 ( .x(n406), .a(n231) );
    inv_1 U304 ( .x(n423), .a(n205) );
    inv_1 U305 ( .x(n426), .a(n199) );
    inv_1 U306 ( .x(n417), .a(n214) );
    inv_1 U307 ( .x(n419), .a(n211) );
    inv_1 U308 ( .x(n420), .a(n208) );
    inv_1 U309 ( .x(n444), .a(n361) );
    inv_1 U310 ( .x(n524), .a(n370) );
    inv_1 U311 ( .x(n450), .a(n356) );
    nand2_1 U312 ( .x(n521), .a(n443), .b(n440) );
    inv_1 U313 ( .x(n372), .a(tc_a[28]) );
    nor2_1 U314 ( .x(n451), .a(n452), .b(n453) );
    nor2_1 U315 ( .x(n458), .a(n459), .b(n460) );
    inv_1 U316 ( .x(n468), .a(n331) );
    nor2_1 U317 ( .x(n464), .a(n465), .b(n466) );
    inv_1 U318 ( .x(n494), .a(n295) );
    nand2_1 U319 ( .x(n273), .a(n274), .b(n275) );
    nand2_1 U320 ( .x(n279), .a(n280), .b(n281) );
    nand2_1 U321 ( .x(n276), .a(n277), .b(n278) );
    nand2_1 U322 ( .x(n262), .a(n263), .b(n264) );
    nand2_1 U323 ( .x(n259), .a(n260), .b(n261) );
    nand2_1 U324 ( .x(n256), .a(n257), .b(n258) );
    nand2_1 U325 ( .x(n253), .a(n254), .b(n255) );
    nand2_1 U326 ( .x(n228), .a(n229), .b(n230) );
    nand2_1 U327 ( .x(n225), .a(n226), .b(n227) );
    nand2_1 U328 ( .x(n219), .a(n220), .b(n221) );
    nand2_1 U329 ( .x(n239), .a(n240), .b(n241) );
    nand2_1 U330 ( .x(n202), .a(n203), .b(n204) );
    nand2_1 U331 ( .x(n196), .a(n197), .b(n198) );
    nor2_1 U332 ( .x(n391), .a(n392), .b(n393) );
    nor2_1 U333 ( .x(n388), .a(n389), .b(n390) );
    nor2_1 U334 ( .x(n381), .a(n382), .b(n126) );
    nor2_1 U335 ( .x(n402), .a(n403), .b(n124) );
    nor2_1 U336 ( .x(n408), .a(n409), .b(n410) );
    inv_1 U337 ( .x(n459), .a(n341) );
    inv_1 U338 ( .x(n465), .a(n328) );
    inv_1 U339 ( .x(n466), .a(n325) );
    inv_1 U340 ( .x(n460), .a(n338) );
    nand2_1 U341 ( .x(n361), .a(n362), .b(n363) );
    nand2_1 U342 ( .x(n373), .a(n374), .b(n375) );
    nand2_1 U343 ( .x(n356), .a(n358), .b(n357) );
    inv_1 U344 ( .x(n452), .a(n352) );
    inv_1 U345 ( .x(n484), .a(n299) );
    inv_1 U346 ( .x(n489), .a(n289) );
    inv_1 U347 ( .x(n492), .a(n286) );
    inv_1 U348 ( .x(n490), .a(n292) );
    inv_1 U349 ( .x(n473), .a(n317) );
    inv_1 U350 ( .x(n471), .a(n322) );
    inv_1 U351 ( .x(n482), .a(n306) );
    inv_1 U352 ( .x(n476), .a(n314) );
    nand2_1 U353 ( .x(n367), .a(n368), .b(n369) );
    nand2_1 U354 ( .x(n331), .a(n332), .b(n333) );
    nand2_1 U355 ( .x(n302), .a(n303), .b(n304) );
    nand2_1 U356 ( .x(n295), .a(n296), .b(n297) );
    inv_1 U357 ( .x(n275), .a(\tc_wd[56] ) );
    inv_1 U358 ( .x(n285), .a(\tc_wd[63] ) );
    inv_1 U359 ( .x(n283), .a(\tc_wd[60] ) );
    inv_1 U360 ( .x(n281), .a(\tc_wd[61] ) );
    inv_1 U361 ( .x(n278), .a(\tc_wd[59] ) );
    inv_1 U362 ( .x(n264), .a(\tc_wd[53] ) );
    inv_1 U363 ( .x(n261), .a(\tc_wd[51] ) );
    inv_1 U364 ( .x(n258), .a(\tc_wd[48] ) );
    inv_1 U365 ( .x(n254), .a(tc_wd[17]) );
    inv_1 U366 ( .x(n255), .a(\tc_wd[49] ) );
    inv_1 U367 ( .x(n230), .a(tc_wd[37]) );
    inv_1 U368 ( .x(n227), .a(tc_wd[35]) );
    inv_1 U369 ( .x(n221), .a(tc_wd[33]) );
    inv_1 U370 ( .x(n241), .a(\tc_wd[40] ) );
    inv_1 U371 ( .x(n204), .a(tc_wd[42]) );
    inv_1 U372 ( .x(n198), .a(tc_wd[34]) );
    nand2_1 U373 ( .x(n341), .a(n342), .b(n343) );
    nand2_1 U374 ( .x(n345), .a(n347), .b(n346) );
    nand2_1 U375 ( .x(n328), .a(n329), .b(n330) );
    nand2_1 U376 ( .x(n325), .a(n326), .b(n327) );
    nand2_1 U377 ( .x(n338), .a(n340), .b(n339) );
    inv_1 U378 ( .x(n362), .a(tc_a[24]) );
    inv_1 U379 ( .x(n363), .a(tc_a[56]) );
    inv_1 U380 ( .x(n357), .a(tc_a[22]) );
    inv_1 U381 ( .x(n358), .a(tc_a[54]) );
    nand2_1 U382 ( .x(n352), .a(n353), .b(n354) );
    nand2_1 U383 ( .x(n299), .a(n300), .b(n301) );
    nand2_1 U384 ( .x(n289), .a(n290), .b(n291) );
    nand2_1 U385 ( .x(n286), .a(n287), .b(n288) );
    nand2_1 U386 ( .x(n292), .a(n293), .b(n294) );
    nand2_1 U387 ( .x(n317), .a(n318), .b(n319) );
    nand2_1 U388 ( .x(n322), .a(n323), .b(n324) );
    nand2_1 U389 ( .x(n306), .a(n307), .b(n308) );
    nand2_1 U390 ( .x(n314), .a(n315), .b(n316) );
    inv_1 U391 ( .x(n332), .a(tc_a[4]) );
    inv_1 U392 ( .x(n333), .a(tc_a[36]) );
    inv_1 U393 ( .x(n296), .a(tc_a[31]) );
    inv_1 U394 ( .x(n342), .a(tc_itag[2]) );
    inv_1 U395 ( .x(n343), .a(tc_itag[7]) );
    inv_1 U396 ( .x(n346), .a(tc_a[15]) );
    inv_1 U397 ( .x(n347), .a(tc_a[47]) );
    inv_1 U398 ( .x(n329), .a(tc_a[2]) );
    inv_1 U399 ( .x(n330), .a(tc_a[34]) );
    inv_1 U400 ( .x(n326), .a(tc_a[5]) );
    inv_1 U401 ( .x(n327), .a(tc_a[37]) );
    inv_1 U402 ( .x(n337), .a(tc_a[62]) );
    inv_1 U403 ( .x(n339), .a(tc_lock[0]) );
    inv_1 U404 ( .x(n340), .a(tc_lock[1]) );
    inv_1 U405 ( .x(n353), .a(tc_a[13]) );
    inv_1 U406 ( .x(n354), .a(tc_a[45]) );
    inv_1 U407 ( .x(n300), .a(tc_a[1]) );
    inv_1 U408 ( .x(n290), .a(tc_a[10]) );
    inv_1 U409 ( .x(n291), .a(tc_a[42]) );
    inv_1 U410 ( .x(n287), .a(tc_seq[0]) );
    inv_1 U411 ( .x(n288), .a(tc_seq[1]) );
    inv_1 U412 ( .x(n293), .a(tc_a[23]) );
    inv_1 U413 ( .x(n294), .a(tc_a[55]) );
    inv_1 U414 ( .x(n318), .a(tc_a[19]) );
    inv_1 U415 ( .x(n323), .a(tc_a[0]) );
    inv_1 U416 ( .x(n307), .a(tc_a[25]) );
    inv_1 U417 ( .x(n308), .a(tc_a[57]) );
    buf_1 U418 ( .x(we_i), .a(tc_rnw[0]) );
    matched_delay_cp2slave_resp_wb U419 ( .x(req_out_delayed), .a(req_out) );
    and4_1 U420 ( .x(_25_net_), .a(sel_o[0]), .b(sel_o[1]), .c(n529), .d(n530)
         );
    inv_1 U421 ( .x(_24_net_), .a(we_i) );
    and2_1 U422 ( .x(tc_defer), .a(rty_o), .b(respond) );
    and4_1 U423 ( .x(_26_net_), .a(sel_o[0]), .b(sel_o[1]), .c(sel_o[3]), .d(
        sel_o[2]) );
    inv_1 U424 ( .x(n532), .a(acc_o) );
    inv_1 U425 ( .x(n531), .a(rty_o) );
    inv_1 U426 ( .x(n529), .a(sel_o[2]) );
    inv_1 U427 ( .x(n530), .a(sel_o[3]) );
    buf_1 U150 ( .x(n142), .a(req_in_i) );
    matched_delay_cp2slave_com_wb matchDelCom ( .x(req_in), .a(req_in_i) );
    nand2_1 U275 ( .x(req_in_i), .a(n186), .b(n187) );
    inv_1 U221 ( .x(n186), .a(all_w) );
    inv_1 U269 ( .x(n187), .a(all_r) );
    dffp_1 mult_i_reg ( .q(mult_i), .d(n137), .ck(n142) );
    ao222_1 \cg_respond/__tmp99/U1  ( .x(respond), .a(req_out), .b(tc_ack), 
        .c(req_out), .d(respond), .e(tc_ack), .f(respond) );
    oa21_1 \cg_all_r/__tmp99/U1  ( .x(all_r), .a(tc_rnw[1]), .b(all_r), .c(
        comp_basic) );
    ao31_1 \cg_all_w/__tmp99/aoi  ( .x(\cg_all_w/__tmp99/loop ), .a(comp_basic
        ), .b(comp_wd), .c(we_i), .d(all_w) );
    oa21_1 \cg_all_w/__tmp99/outGate  ( .x(all_w), .a(comp_basic), .b(comp_wd), 
        .c(\cg_all_w/__tmp99/loop ) );
    ao222_1 \cg_wd/__tmp99/U1  ( .x(comp_wd), .a(complw0), .b(complw1), .c(
        complw0), .d(comp_wd), .e(complw1), .f(comp_wd) );
    ao222_1 \cg_basic/__tmp99/U1  ( .x(comp_basic), .a(complb0), .b(complb1), 
        .c(complb0), .d(comp_basic), .e(complb1), .f(comp_basic) );
    inv_1 \Usze1/Uii  ( .x(\Usze1/ni ), .a(_26_net_) );
    inv_1 \Usze1/Uih  ( .x(\Usze1/nh ), .a(tr_size[3]) );
    inv_1 \Usze1/Uil  ( .x(\Usze1/nl ), .a(tr_size[1]) );
    ao23_1 \Usze1/Ucl/U1/U1  ( .x(tr_size[1]), .a(n2), .b(tr_size[1]), .c(n1), 
        .d(\Usze1/ni ), .e(\Usze1/nh ) );
    ao23_1 \Usze1/Uch/U1/U1  ( .x(tr_size[3]), .a(n1), .b(tr_size[3]), .c(n1), 
        .d(_26_net_), .e(\Usze1/nl ) );
    inv_1 \Usze0/Uii  ( .x(\Usze0/ni ), .a(_25_net_) );
    inv_1 \Usze0/Uih  ( .x(\Usze0/nh ), .a(tr_size[2]) );
    inv_1 \Usze0/Uil  ( .x(\Usze0/nl ), .a(tr_size[0]) );
    ao23_1 \Usze0/Ucl/U1/U1  ( .x(tr_size[0]), .a(n2), .b(tr_size[0]), .c(n1), 
        .d(\Usze0/ni ), .e(\Usze0/nh ) );
    ao23_1 \Usze0/Uch/U1/U1  ( .x(tr_size[2]), .a(n2), .b(tr_size[2]), .c(n1), 
        .d(_25_net_), .e(\Usze0/nl ) );
    inv_1 \Urnw/Uii  ( .x(\Urnw/ni ), .a(_24_net_) );
    inv_1 \Urnw/Uih  ( .x(\Urnw/nh ), .a(tr_rnw[1]) );
    inv_1 \Urnw/Uil  ( .x(\Urnw/nl ), .a(tr_rnw[0]) );
    ao23_1 \Urnw/Ucl/U1/U1  ( .x(tr_rnw[0]), .a(n1), .b(tr_rnw[0]), .c(n1), 
        .d(\Urnw/ni ), .e(\Urnw/nh ) );
    ao23_1 \Urnw/Uch/U1/U1  ( .x(tr_rnw[1]), .a(n1), .b(tr_rnw[1]), .c(n1), 
        .d(_24_net_), .e(\Urnw/nl ) );
    inv_1 \Uerr/Uii  ( .x(\Uerr/ni ), .a(err_o) );
    inv_1 \Uerr/Uih  ( .x(\Uerr/nh ), .a(tr_err[1]) );
    inv_1 \Uerr/Uil  ( .x(\Uerr/nl ), .a(tr_err[0]) );
    ao23_1 \Uerr/Ucl/U1/U1  ( .x(tr_err[0]), .a(n1), .b(tr_err[0]), .c(n1), 
        .d(\Uerr/ni ), .e(\Uerr/nh ) );
    ao23_1 \Uerr/Uch/U1/U1  ( .x(tr_err[1]), .a(n1), .b(tr_err[1]), .c(n1), 
        .d(err_o), .e(\Uerr/nl ) );
    inv_0 U1 ( .x(n298), .a(tc_itag[6]) );
    nor2_0 U2 ( .x(n485), .a(tc_itag[1]), .b(tc_itag[6]) );
    inv_0 U4 ( .x(n344), .a(tc_itag[8]) );
    nor2_0 U8 ( .x(n462), .a(tc_itag[3]), .b(tc_itag[8]) );
    nor2_0 U92 ( .x(n496), .a(tc_size[0]), .b(tc_size[1]) );
    nor2_0 U93 ( .x(n194), .a(tc_size[0]), .b(tc_size[2]) );
    buf_16 U104 ( .x(n1), .a(req_out_delayed) );
    buf_16 U111 ( .x(n2), .a(req_out_delayed) );
endmodule


module slave_if_wb ( nReset, sc_req, sc_we, sc_mult, sc_seq, sc_prd, sc_ts, 
    sc_st, sc_sel, sc_adr, sc_dat, sc_ack, sr_req, sr_err, sr_rty, sr_acc, 
    sr_mult, sr_ts, sr_rt, sr_sel, sr_dat, sr_ack, chaincommand, 
    nchaincommandack, chainresponse, nchainresponseack, e_dp, e_ip, e_tic, 
    r_dp, r_ip, r_tic );
output [2:0] sc_ts;
output [4:0] sc_st;
output [3:0] sc_sel;
output [31:0] sc_adr;
output [31:0] sc_dat;
input  [2:0] sr_ts;
input  [4:0] sr_rt;
input  [3:0] sr_sel;
input  [31:0] sr_dat;
input  [4:0] chaincommand;
output [4:0] chainresponse;
input  [2:0] e_dp;
input  [2:0] e_ip;
input  [2:0] e_tic;
input  [2:0] r_dp;
input  [2:0] r_ip;
input  [2:0] r_tic;
input  nReset, sc_ack, sr_req, sr_err, sr_rty, sr_acc, sr_mult, 
    nchainresponseack;
output sc_req, sc_we, sc_mult, sc_seq, sc_prd, sr_ack, nchaincommandack;
    wire \ct_a[63] , \ct_a[62] , \ct_a[61] , \ct_a[60] , \ct_a[59] , 
        \ct_a[58] , \ct_a[57] , \ct_a[56] , \ct_a[55] , \ct_a[54] , \ct_a[53] , 
        \ct_a[52] , \ct_a[51] , \ct_a[50] , \ct_a[49] , \ct_a[48] , \ct_a[47] , 
        \ct_a[46] , \ct_a[45] , \ct_a[44] , \ct_a[43] , \ct_a[42] , \ct_a[41] , 
        \ct_a[40] , \ct_a[39] , \ct_a[38] , \ct_a[37] , \ct_a[36] , \ct_a[35] , 
        \ct_a[34] , \ct_a[33] , \ct_a[32] , \ct_a[31] , \ct_a[30] , \ct_a[29] , 
        \ct_a[28] , \ct_a[27] , \ct_a[26] , \ct_a[25] , \ct_a[24] , \ct_a[23] , 
        \ct_a[22] , \ct_a[21] , \ct_a[20] , \ct_a[19] , \ct_a[18] , \ct_a[17] , 
        \ct_a[16] , \ct_a[15] , \ct_a[14] , \ct_a[13] , \ct_a[12] , \ct_a[11] , 
        \ct_a[10] , \ct_a[9] , \ct_a[8] , \ct_a[7] , \ct_a[6] , \ct_a[5] , 
        \ct_a[4] , \ct_a[3] , \ct_a[2] , \ct_a[1] , \ct_a[0] , \ct_wd[63] , 
        \ct_wd[62] , \ct_wd[61] , \ct_wd[60] , \ct_wd[59] , \ct_wd[58] , 
        \ct_wd[57] , \ct_wd[56] , \ct_wd[55] , \ct_wd[54] , \ct_wd[53] , 
        \ct_wd[52] , \ct_wd[51] , \ct_wd[50] , \ct_wd[49] , \ct_wd[48] , 
        \ct_wd[47] , \ct_wd[46] , \ct_wd[45] , \ct_wd[44] , \ct_wd[43] , 
        \ct_wd[42] , \ct_wd[41] , \ct_wd[40] , \ct_wd[39] , \ct_wd[38] , 
        \ct_wd[37] , \ct_wd[36] , \ct_wd[35] , \ct_wd[34] , \ct_wd[33] , 
        \ct_wd[32] , \ct_wd[31] , \ct_wd[30] , \ct_wd[29] , \ct_wd[28] , 
        \ct_wd[27] , \ct_wd[26] , \ct_wd[25] , \ct_wd[24] , \ct_wd[23] , 
        \ct_wd[22] , \ct_wd[21] , \ct_wd[20] , \ct_wd[19] , \ct_wd[18] , 
        \ct_wd[17] , \ct_wd[16] , \ct_wd[15] , \ct_wd[14] , \ct_wd[13] , 
        \ct_wd[12] , \ct_wd[11] , \ct_wd[10] , \ct_wd[9] , \ct_wd[8] , 
        \ct_wd[7] , \ct_wd[6] , \ct_wd[5] , \ct_wd[4] , \ct_wd[3] , \ct_wd[2] , 
        \ct_wd[1] , \ct_wd[0] , \ct_rnw[1] , \ct_rnw[0] , \ct_lock[1] , 
        \ct_lock[0] , \ct_seq[1] , \ct_seq[0] , \ct_size[3] , \ct_size[2] , 
        \ct_size[1] , \ct_size[0] , \ct_itag[9] , \ct_itag[8] , \ct_itag[7] , 
        \ct_itag[6] , \ct_itag[5] , \ct_itag[4] , \ct_itag[3] , \ct_itag[2] , 
        \ct_itag[1] , \ct_itag[0] , ct_ack, ct_ok, ct_defer, ct_slow, 
        \rt_rd[63] , \rt_rd[62] , \rt_rd[61] , \rt_rd[60] , \rt_rd[59] , 
        \rt_rd[58] , \rt_rd[57] , \rt_rd[56] , \rt_rd[55] , \rt_rd[54] , 
        \rt_rd[53] , \rt_rd[52] , \rt_rd[51] , \rt_rd[50] , \rt_rd[49] , 
        \rt_rd[48] , \rt_rd[47] , \rt_rd[46] , \rt_rd[45] , \rt_rd[44] , 
        \rt_rd[43] , \rt_rd[42] , \rt_rd[41] , \rt_rd[40] , \rt_rd[39] , 
        \rt_rd[38] , \rt_rd[37] , \rt_rd[36] , \rt_rd[35] , \rt_rd[34] , 
        \rt_rd[33] , \rt_rd[32] , \rt_rd[31] , \rt_rd[30] , \rt_rd[29] , 
        \rt_rd[28] , \rt_rd[27] , \rt_rd[26] , \rt_rd[25] , \rt_rd[24] , 
        \rt_rd[23] , \rt_rd[22] , \rt_rd[21] , \rt_rd[20] , \rt_rd[19] , 
        \rt_rd[18] , \rt_rd[17] , \rt_rd[16] , \rt_rd[15] , \rt_rd[14] , 
        \rt_rd[13] , \rt_rd[12] , \rt_rd[11] , \rt_rd[10] , \rt_rd[9] , 
        \rt_rd[8] , \rt_rd[7] , \rt_rd[6] , \rt_rd[5] , \rt_rd[4] , \rt_rd[3] , 
        \rt_rd[2] , \rt_rd[1] , \rt_rd[0] , \rt_err[1] , \rt_err[0] , rt_ack, 
        \tag_h[4] , \tag_h[3] , \tag_h[2] , \tag_h[1] , \tag_h[0] , \tag_l[4] , 
        \tag_l[3] , \tag_l[2] , \tag_l[1] , \tag_l[0] , \route[4] , \route[1] , 
        \route[0] , nroute_ack, routetx_req, routetx_ack, \eh[1] , \eh[0] , 
        \el[2] , \el[1] , \el[0] , \rh[2] , \rh[1] , \rl[2] , \rl[1] , \rl[0] , 
        reset;
    wire SYNOPSYS_UNCONNECTED_1 , SYNOPSYS_UNCONNECTED_2 , 
	SYNOPSYS_UNCONNECTED_3 , SYNOPSYS_UNCONNECTED_4 , SYNOPSYS_UNCONNECTED_5 ;
    assign sc_prd = 1'b0;
    assign sc_ts[2] = 1'b0;
    assign sc_ts[1] = 1'b0;
    assign sc_ts[0] = 1'b0;
    assign sc_sel[0] = 1'b1;
    target_wb tg ( .addr({\ct_a[63] , \ct_a[62] , \ct_a[61] , \ct_a[60] , 
        \ct_a[59] , \ct_a[58] , \ct_a[57] , \ct_a[56] , \ct_a[55] , \ct_a[54] , 
        \ct_a[53] , \ct_a[52] , \ct_a[51] , \ct_a[50] , \ct_a[49] , \ct_a[48] , 
        \ct_a[47] , \ct_a[46] , \ct_a[45] , \ct_a[44] , \ct_a[43] , \ct_a[42] , 
        \ct_a[41] , \ct_a[40] , \ct_a[39] , \ct_a[38] , \ct_a[37] , \ct_a[36] , 
        \ct_a[35] , \ct_a[34] , \ct_a[33] , \ct_a[32] , \ct_a[31] , \ct_a[30] , 
        \ct_a[29] , \ct_a[28] , \ct_a[27] , \ct_a[26] , \ct_a[25] , \ct_a[24] , 
        \ct_a[23] , \ct_a[22] , \ct_a[21] , \ct_a[20] , \ct_a[19] , \ct_a[18] , 
        \ct_a[17] , \ct_a[16] , \ct_a[15] , \ct_a[14] , \ct_a[13] , \ct_a[12] , 
        \ct_a[11] , \ct_a[10] , \ct_a[9] , \ct_a[8] , \ct_a[7] , \ct_a[6] , 
        \ct_a[5] , \ct_a[4] , \ct_a[3] , \ct_a[2] , \ct_a[1] , \ct_a[0] }), 
        .chainresponse(chainresponse), .crnw({\ct_rnw[1] , \ct_rnw[0] }), 
        .csize({\ct_size[3] , \ct_size[2] , \ct_size[1] , \ct_size[0] }), 
        .ctag({\ct_itag[9] , \ct_itag[8] , \ct_itag[7] , \ct_itag[6] , 
        \ct_itag[5] , \ct_itag[4] , \ct_itag[3] , \ct_itag[2] , \ct_itag[1] , 
        \ct_itag[0] }), .lock({\ct_lock[1] , \ct_lock[0] }), 
        .nchaincommandack(nchaincommandack), .nrouteack(nroute_ack), .rack(
        rt_ack), .routetxreq(routetx_req), .seq({\ct_seq[1] , \ct_seq[0] }), 
        .tag_h({\tag_h[4] , \tag_h[3] , \tag_h[2] , \tag_h[1] , \tag_h[0] }), 
        .tag_l({\tag_l[4] , \tag_l[3] , \tag_l[2] , \tag_l[1] , \tag_l[0] }), 
        .wd({\ct_wd[63] , \ct_wd[62] , \ct_wd[61] , \ct_wd[60] , \ct_wd[59] , 
        \ct_wd[58] , \ct_wd[57] , \ct_wd[56] , \ct_wd[55] , \ct_wd[54] , 
        \ct_wd[53] , \ct_wd[52] , \ct_wd[51] , \ct_wd[50] , \ct_wd[49] , 
        \ct_wd[48] , \ct_wd[47] , \ct_wd[46] , \ct_wd[45] , \ct_wd[44] , 
        \ct_wd[43] , \ct_wd[42] , \ct_wd[41] , \ct_wd[40] , \ct_wd[39] , 
        \ct_wd[38] , \ct_wd[37] , \ct_wd[36] , \ct_wd[35] , \ct_wd[34] , 
        \ct_wd[33] , \ct_wd[32] , \ct_wd[31] , \ct_wd[30] , \ct_wd[29] , 
        \ct_wd[28] , \ct_wd[27] , \ct_wd[26] , \ct_wd[25] , \ct_wd[24] , 
        \ct_wd[23] , \ct_wd[22] , \ct_wd[21] , \ct_wd[20] , \ct_wd[19] , 
        \ct_wd[18] , \ct_wd[17] , \ct_wd[16] , \ct_wd[15] , \ct_wd[14] , 
        \ct_wd[13] , \ct_wd[12] , \ct_wd[11] , \ct_wd[10] , \ct_wd[9] , 
        \ct_wd[8] , \ct_wd[7] , \ct_wd[6] , \ct_wd[5] , \ct_wd[4] , \ct_wd[3] , 
        \ct_wd[2] , \ct_wd[1] , \ct_wd[0] }), .cack(ct_ack), .cdefer(ct_defer), 
        .chaincommand(chaincommand), .cndefer(ct_slow), .cok(ct_ok), .err({
        \rt_err[1] , \rt_err[0] }), .nReset(nReset), .nchainresponseack(
        nchainresponseack), .rd({\rt_rd[63] , \rt_rd[62] , \rt_rd[61] , 
        \rt_rd[60] , \rt_rd[59] , \rt_rd[58] , \rt_rd[57] , \rt_rd[56] , 
        \rt_rd[55] , \rt_rd[54] , \rt_rd[53] , \rt_rd[52] , \rt_rd[51] , 
        \rt_rd[50] , \rt_rd[49] , \rt_rd[48] , \rt_rd[47] , \rt_rd[46] , 
        \rt_rd[45] , \rt_rd[44] , \rt_rd[43] , \rt_rd[42] , \rt_rd[41] , 
        \rt_rd[40] , \rt_rd[39] , \rt_rd[38] , \rt_rd[37] , \rt_rd[36] , 
        \rt_rd[35] , \rt_rd[34] , \rt_rd[33] , \rt_rd[32] , \rt_rd[31] , 
        \rt_rd[30] , \rt_rd[29] , \rt_rd[28] , \rt_rd[27] , \rt_rd[26] , 
        \rt_rd[25] , \rt_rd[24] , \rt_rd[23] , \rt_rd[22] , \rt_rd[21] , 
        \rt_rd[20] , \rt_rd[19] , \rt_rd[18] , \rt_rd[17] , \rt_rd[16] , 
        \rt_rd[15] , \rt_rd[14] , \rt_rd[13] , \rt_rd[12] , \rt_rd[11] , 
        \rt_rd[10] , \rt_rd[9] , \rt_rd[8] , \rt_rd[7] , \rt_rd[6] , 
        \rt_rd[5] , \rt_rd[4] , \rt_rd[3] , \rt_rd[2] , \rt_rd[1] , \rt_rd[0] 
        }), .route({\route[4] , 1'b0, 1'b0, \route[1] , \route[0] }), 
        .routetxack(routetx_ack) );
    t_adec_wb dec ( .e_h({SYNOPSYS_UNCONNECTED_1, \eh[1] , \eh[0] }), .e_l({
        \el[2] , \el[1] , \el[0] }), .r_h({\rh[2] , \rh[1] , 
        SYNOPSYS_UNCONNECTED_2}), .r_l({\rl[2] , \rl[1] , \rl[0] }), .e_dp(
        e_dp), .e_ip(e_ip), .e_tic(e_tic), .r_dp(r_dp), .r_ip(r_ip), .r_tic(
        r_tic), .tag_h({\tag_h[4] , \tag_h[3] , \tag_h[2] , \tag_h[1] , 
        \tag_h[0] }), .tag_l({\tag_l[4] , \tag_l[3] , \tag_l[2] , \tag_l[1] , 
        \tag_l[0] }) );
    resp_route_tx_wb rt ( .o({\route[4] , SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, \route[1] , \route[0] }), .rtxack(routetx_ack), 
        .e_h({1'b0, \eh[1] , \eh[0] }), .e_l({\el[2] , \el[1] , \el[0] }), 
        .noa(nroute_ack), .r_h({\rh[2] , \rh[1] , 1'b0}), .r_l({\rl[2] , 
        \rl[1] , \rl[0] }), .rtxreq(routetx_req) );
    inv_2 U1 ( .x(reset), .a(nReset) );
    cp2slave_wb chainif2slave ( .tc_seq({\ct_seq[1] , \ct_seq[0] }), .tc_size(
        {\ct_size[3] , \ct_size[2] , \ct_size[1] , \ct_size[0] }), .tc_itag({
        \ct_itag[9] , \ct_itag[8] , \ct_itag[7] , \ct_itag[6] , \ct_itag[5] , 
        \ct_itag[4] , \ct_itag[3] , \ct_itag[2] , \ct_itag[1] , \ct_itag[0] }), 
        .tc_wd({\ct_wd[63] , \ct_wd[62] , \ct_wd[61] , \ct_wd[60] , 
        \ct_wd[59] , \ct_wd[58] , \ct_wd[57] , \ct_wd[56] , \ct_wd[55] , 
        \ct_wd[54] , \ct_wd[53] , \ct_wd[52] , \ct_wd[51] , \ct_wd[50] , 
        \ct_wd[49] , \ct_wd[48] , \ct_wd[47] , \ct_wd[46] , \ct_wd[45] , 
        \ct_wd[44] , \ct_wd[43] , \ct_wd[42] , \ct_wd[41] , \ct_wd[40] , 
        \ct_wd[39] , \ct_wd[38] , \ct_wd[37] , \ct_wd[36] , \ct_wd[35] , 
        \ct_wd[34] , \ct_wd[33] , \ct_wd[32] , \ct_wd[31] , \ct_wd[30] , 
        \ct_wd[29] , \ct_wd[28] , \ct_wd[27] , \ct_wd[26] , \ct_wd[25] , 
        \ct_wd[24] , \ct_wd[23] , \ct_wd[22] , \ct_wd[21] , \ct_wd[20] , 
        \ct_wd[19] , \ct_wd[18] , \ct_wd[17] , \ct_wd[16] , \ct_wd[15] , 
        \ct_wd[14] , \ct_wd[13] , \ct_wd[12] , \ct_wd[11] , \ct_wd[10] , 
        \ct_wd[9] , \ct_wd[8] , \ct_wd[7] , \ct_wd[6] , \ct_wd[5] , \ct_wd[4] , 
        \ct_wd[3] , \ct_wd[2] , \ct_wd[1] , \ct_wd[0] }), .tc_lock({
        \ct_lock[1] , \ct_lock[0] }), .tc_a({\ct_a[63] , \ct_a[62] , 
        \ct_a[61] , \ct_a[60] , \ct_a[59] , \ct_a[58] , \ct_a[57] , \ct_a[56] , 
        \ct_a[55] , \ct_a[54] , \ct_a[53] , \ct_a[52] , \ct_a[51] , \ct_a[50] , 
        \ct_a[49] , \ct_a[48] , \ct_a[47] , \ct_a[46] , \ct_a[45] , \ct_a[44] , 
        \ct_a[43] , \ct_a[42] , \ct_a[41] , \ct_a[40] , \ct_a[39] , \ct_a[38] , 
        \ct_a[37] , \ct_a[36] , \ct_a[35] , \ct_a[34] , \ct_a[33] , \ct_a[32] , 
        \ct_a[31] , \ct_a[30] , \ct_a[29] , \ct_a[28] , \ct_a[27] , \ct_a[26] , 
        \ct_a[25] , \ct_a[24] , \ct_a[23] , \ct_a[22] , \ct_a[21] , \ct_a[20] , 
        \ct_a[19] , \ct_a[18] , \ct_a[17] , \ct_a[16] , \ct_a[15] , \ct_a[14] , 
        \ct_a[13] , \ct_a[12] , \ct_a[11] , \ct_a[10] , \ct_a[9] , \ct_a[8] , 
        \ct_a[7] , \ct_a[6] , \ct_a[5] , \ct_a[4] , \ct_a[3] , \ct_a[2] , 
        \ct_a[1] , \ct_a[0] }), .tc_rnw({\ct_rnw[1] , \ct_rnw[0] }), .tc_ok(
        ct_ok), .tc_defer(ct_defer), .tc_slow(ct_slow), .tc_ack(ct_ack), 
        .req_in(sc_req), .st_i(sc_st), .we_i(sc_we), .mult_i(sc_mult), .adr_i(
        sc_adr), .dat_i(sc_dat), .seq_i(sc_seq), .sel_i({sc_sel[3], sc_sel[2], 
        sc_sel[1], SYNOPSYS_UNCONNECTED_5}), .ack_in(sc_ack), .tr_rd({
        \rt_rd[63] , \rt_rd[62] , \rt_rd[61] , \rt_rd[60] , \rt_rd[59] , 
        \rt_rd[58] , \rt_rd[57] , \rt_rd[56] , \rt_rd[55] , \rt_rd[54] , 
        \rt_rd[53] , \rt_rd[52] , \rt_rd[51] , \rt_rd[50] , \rt_rd[49] , 
        \rt_rd[48] , \rt_rd[47] , \rt_rd[46] , \rt_rd[45] , \rt_rd[44] , 
        \rt_rd[43] , \rt_rd[42] , \rt_rd[41] , \rt_rd[40] , \rt_rd[39] , 
        \rt_rd[38] , \rt_rd[37] , \rt_rd[36] , \rt_rd[35] , \rt_rd[34] , 
        \rt_rd[33] , \rt_rd[32] , \rt_rd[31] , \rt_rd[30] , \rt_rd[29] , 
        \rt_rd[28] , \rt_rd[27] , \rt_rd[26] , \rt_rd[25] , \rt_rd[24] , 
        \rt_rd[23] , \rt_rd[22] , \rt_rd[21] , \rt_rd[20] , \rt_rd[19] , 
        \rt_rd[18] , \rt_rd[17] , \rt_rd[16] , \rt_rd[15] , \rt_rd[14] , 
        \rt_rd[13] , \rt_rd[12] , \rt_rd[11] , \rt_rd[10] , \rt_rd[9] , 
        \rt_rd[8] , \rt_rd[7] , \rt_rd[6] , \rt_rd[5] , \rt_rd[4] , \rt_rd[3] , 
        \rt_rd[2] , \rt_rd[1] , \rt_rd[0] }), .tr_err({\rt_err[1] , 
        \rt_err[0] }), .tr_ack(rt_ack), .req_out(sr_req), .dat_o(sr_dat), 
        .err_o(sr_err), .rty_o(sr_rty), .acc_o(sr_acc), .sel_o(sr_sel), 
        .mult_o(sr_mult), .rt_o(sr_rt), .ack_out(sr_ack), .reset(reset) );
endmodule


module wb_block ( nReset, clk, chaincommand, nchaincommandack, chainresponse, 
    nchainresponseack, e_dp, e_ip, e_tic, r_dp, r_ip, r_tic, wb_we_o, 
    wb_stb_cyc_o, wb_ack_i, wb_adr_o, wb_dat_i, wb_dat_o );
input  [4:0] chaincommand;
output [4:0] chainresponse;
input  [2:0] e_dp;
input  [2:0] e_ip;
input  [2:0] e_tic;
input  [2:0] r_dp;
input  [2:0] r_ip;
input  [2:0] r_tic;
output [11:0] wb_adr_o;
input  [31:0] wb_dat_i;
output [31:0] wb_dat_o;
input  nReset, clk, nchainresponseack, wb_ack_i;
output nchaincommandack, wb_we_o, wb_stb_cyc_o;
    wire \sc_st[4] , \sc_st[3] , \sc_st[2] , \sc_st[1] , \sc_st[0] , sc_req, 
        sc_we, \sc_adr[13] , \sc_adr[12] , \sc_adr[11] , \sc_adr[10] , 
        \sc_adr[9] , \sc_adr[8] , \sc_adr[7] , \sc_adr[6] , \sc_adr[5] , 
        \sc_adr[4] , \sc_adr[3] , \sc_adr[2] , \sc_dat[31] , \sc_dat[30] , 
        \sc_dat[29] , \sc_dat[28] , \sc_dat[27] , \sc_dat[26] , \sc_dat[25] , 
        \sc_dat[24] , \sc_dat[23] , \sc_dat[22] , \sc_dat[21] , \sc_dat[20] , 
        \sc_dat[19] , \sc_dat[18] , \sc_dat[17] , \sc_dat[16] , \sc_dat[15] , 
        \sc_dat[14] , \sc_dat[13] , \sc_dat[12] , \sc_dat[11] , \sc_dat[10] , 
        \sc_dat[9] , \sc_dat[8] , \sc_dat[7] , \sc_dat[6] , \sc_dat[5] , 
        \sc_dat[4] , \sc_dat[3] , \sc_dat[2] , \sc_dat[1] , \sc_dat[0] , 
        sc_ack, sr_req, \sr_dat[31] , \sr_dat[30] , \sr_dat[29] , \sr_dat[28] , 
        \sr_dat[27] , \sr_dat[26] , \sr_dat[25] , \sr_dat[24] , \sr_dat[23] , 
        \sr_dat[22] , \sr_dat[21] , \sr_dat[20] , \sr_dat[19] , \sr_dat[18] , 
        \sr_dat[17] , \sr_dat[16] , \sr_dat[15] , \sr_dat[14] , \sr_dat[13] , 
        \sr_dat[12] , \sr_dat[11] , \sr_dat[10] , \sr_dat[9] , \sr_dat[8] , 
        \sr_dat[7] , \sr_dat[6] , \sr_dat[5] , \sr_dat[4] , \sr_dat[3] , 
        \sr_dat[2] , \sr_dat[1] , \sr_dat[0] , sr_ack;
    wire SYNOPSYS_UNCONNECTED_1 , SYNOPSYS_UNCONNECTED_2 , 
	SYNOPSYS_UNCONNECTED_3 , SYNOPSYS_UNCONNECTED_4 , SYNOPSYS_UNCONNECTED_5 , 
	SYNOPSYS_UNCONNECTED_6 , SYNOPSYS_UNCONNECTED_7 , SYNOPSYS_UNCONNECTED_8 , 
	SYNOPSYS_UNCONNECTED_9 , SYNOPSYS_UNCONNECTED_10 , SYNOPSYS_UNCONNECTED_11 , 
	SYNOPSYS_UNCONNECTED_12 , SYNOPSYS_UNCONNECTED_13 , SYNOPSYS_UNCONNECTED_14 , 
	SYNOPSYS_UNCONNECTED_15 , SYNOPSYS_UNCONNECTED_16 , SYNOPSYS_UNCONNECTED_17 , 
	SYNOPSYS_UNCONNECTED_18 , SYNOPSYS_UNCONNECTED_19 , SYNOPSYS_UNCONNECTED_20 ;
    slave_if_wb wbIf ( .nReset(nReset), .sc_req(sc_req), .sc_we(sc_we), 
        .sc_st({\sc_st[4] , \sc_st[3] , \sc_st[2] , \sc_st[1] , \sc_st[0] }), 
        .sc_adr({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, \sc_adr[13] , 
        \sc_adr[12] , \sc_adr[11] , \sc_adr[10] , \sc_adr[9] , \sc_adr[8] , 
        \sc_adr[7] , \sc_adr[6] , \sc_adr[5] , \sc_adr[4] , \sc_adr[3] , 
        \sc_adr[2] , SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20}), 
        .sc_dat({\sc_dat[31] , \sc_dat[30] , \sc_dat[29] , \sc_dat[28] , 
        \sc_dat[27] , \sc_dat[26] , \sc_dat[25] , \sc_dat[24] , \sc_dat[23] , 
        \sc_dat[22] , \sc_dat[21] , \sc_dat[20] , \sc_dat[19] , \sc_dat[18] , 
        \sc_dat[17] , \sc_dat[16] , \sc_dat[15] , \sc_dat[14] , \sc_dat[13] , 
        \sc_dat[12] , \sc_dat[11] , \sc_dat[10] , \sc_dat[9] , \sc_dat[8] , 
        \sc_dat[7] , \sc_dat[6] , \sc_dat[5] , \sc_dat[4] , \sc_dat[3] , 
        \sc_dat[2] , \sc_dat[1] , \sc_dat[0] }), .sc_ack(sc_ack), .sr_req(
        sr_req), .sr_err(1'b0), .sr_rty(1'b0), .sr_acc(1'b0), .sr_mult(1'b0), 
        .sr_ts({1'b0, 1'b0, 1'b0}), .sr_rt({\sc_st[4] , \sc_st[3] , \sc_st[2] , 
        \sc_st[1] , \sc_st[0] }), .sr_sel({1'b1, 1'b1, 1'b1, 1'b1}), .sr_dat({
        \sr_dat[31] , \sr_dat[30] , \sr_dat[29] , \sr_dat[28] , \sr_dat[27] , 
        \sr_dat[26] , \sr_dat[25] , \sr_dat[24] , \sr_dat[23] , \sr_dat[22] , 
        \sr_dat[21] , \sr_dat[20] , \sr_dat[19] , \sr_dat[18] , \sr_dat[17] , 
        \sr_dat[16] , \sr_dat[15] , \sr_dat[14] , \sr_dat[13] , \sr_dat[12] , 
        \sr_dat[11] , \sr_dat[10] , \sr_dat[9] , \sr_dat[8] , \sr_dat[7] , 
        \sr_dat[6] , \sr_dat[5] , \sr_dat[4] , \sr_dat[3] , \sr_dat[2] , 
        \sr_dat[1] , \sr_dat[0] }), .sr_ack(sr_ack), .chaincommand(
        chaincommand), .nchaincommandack(nchaincommandack), .chainresponse(
        chainresponse), .nchainresponseack(nchainresponseack), .e_dp(e_dp), 
        .e_ip(e_ip), .e_tic(e_tic), .r_dp(r_dp), .r_ip(r_ip), .r_tic(r_tic) );
    wishbone wbconv ( .reset_b(nReset), .clk(clk), .ch_we_i(sc_we), .ch_dat_i(
        {\sc_dat[31] , \sc_dat[30] , \sc_dat[29] , \sc_dat[28] , \sc_dat[27] , 
        \sc_dat[26] , \sc_dat[25] , \sc_dat[24] , \sc_dat[23] , \sc_dat[22] , 
        \sc_dat[21] , \sc_dat[20] , \sc_dat[19] , \sc_dat[18] , \sc_dat[17] , 
        \sc_dat[16] , \sc_dat[15] , \sc_dat[14] , \sc_dat[13] , \sc_dat[12] , 
        \sc_dat[11] , \sc_dat[10] , \sc_dat[9] , \sc_dat[8] , \sc_dat[7] , 
        \sc_dat[6] , \sc_dat[5] , \sc_dat[4] , \sc_dat[3] , \sc_dat[2] , 
        \sc_dat[1] , \sc_dat[0] }), .ch_adr_i({\sc_adr[13] , \sc_adr[12] , 
        \sc_adr[11] , \sc_adr[10] , \sc_adr[9] , \sc_adr[8] , \sc_adr[7] , 
        \sc_adr[6] , \sc_adr[5] , \sc_adr[4] , \sc_adr[3] , \sc_adr[2] }), 
        .ch_req_i(sc_req), .ch_ack_i(sc_ack), .ch_req_o(sr_req), .ch_dat_o({
        \sr_dat[31] , \sr_dat[30] , \sr_dat[29] , \sr_dat[28] , \sr_dat[27] , 
        \sr_dat[26] , \sr_dat[25] , \sr_dat[24] , \sr_dat[23] , \sr_dat[22] , 
        \sr_dat[21] , \sr_dat[20] , \sr_dat[19] , \sr_dat[18] , \sr_dat[17] , 
        \sr_dat[16] , \sr_dat[15] , \sr_dat[14] , \sr_dat[13] , \sr_dat[12] , 
        \sr_dat[11] , \sr_dat[10] , \sr_dat[9] , \sr_dat[8] , \sr_dat[7] , 
        \sr_dat[6] , \sr_dat[5] , \sr_dat[4] , \sr_dat[3] , \sr_dat[2] , 
        \sr_dat[1] , \sr_dat[0] }), .ch_ack_o(sr_ack), .wb_we_o(wb_we_o), 
        .wb_stb_cyc_o(wb_stb_cyc_o), .wb_dat_o(wb_dat_o), .wb_adr_o(wb_adr_o), 
        .wb_dat_i(wb_dat_i), .wb_ack_i(wb_ack_i) );
endmodule


module i_adec_iport ( e_h, e_l, r_h, r_l, ah, al, e_bare, e_dm, e_im, e_wish, 
    r_bare, r_dm, r_im, r_wish, force_bare );
output [3:0] e_h;
output [3:0] e_l;
output [3:0] r_h;
output [3:0] r_l;
input  [31:0] ah;
input  [31:0] al;
input  [3:0] e_bare;
input  [3:0] e_dm;
input  [3:0] e_im;
input  [3:0] e_wish;
input  [3:0] r_bare;
input  [3:0] r_dm;
input  [3:0] r_im;
input  [3:0] r_wish;
input  force_bare;
    wire \e_l[2] , \e_h[0] , n14, n15, \r_l[2] , \r_l[0] , im_i, dm_i, wish_i, 
        bare_i, n1, n2, n3, n6, n7, \e_l[3] , \e_l[0] , n12;
    assign e_h[3] = 1'b0;
    assign e_h[0] = \e_h[0] ;
    assign e_l[3] = \e_l[3] ;
    assign e_l[2] = \e_l[2] ;
    assign e_l[0] = \e_l[0] ;
    assign r_h[3] = \e_l[2] ;
    assign r_h[2] = \e_h[0] ;
    assign r_h[0] = 1'b0;
    assign r_l[2] = \e_l[0] ;
    assign r_l[0] = \e_l[3] ;
    ao222_1 \U1632/U18/U1/U1  ( .x(wish_i), .a(n6), .b(al[30]), .c(n6), .d(
        wish_i), .e(al[30]), .f(wish_i) );
    ao222_1 \U1633/U18/U1/U1  ( .x(bare_i), .a(n6), .b(ah[30]), .c(n6), .d(
        bare_i), .e(ah[30]), .f(bare_i) );
    ao222_1 \U1634/U18/U1/U1  ( .x(im_i), .a(al[11]), .b(n7), .c(al[11]), .d(
        im_i), .e(n7), .f(im_i) );
    ao222_1 \U1635/U18/U1/U1  ( .x(dm_i), .a(ah[11]), .b(n7), .c(ah[11]), .d(
        dm_i), .e(n7), .f(dm_i) );
    or3_1 U1 ( .x(\r_l[2] ), .a(wish_i), .b(bare_i), .c(force_bare) );
    or2_1 U2 ( .x(r_l[1]), .a(\e_l[0] ), .b(im_i) );
    or2_1 U3 ( .x(\r_l[0] ), .a(dm_i), .b(r_l[1]) );
    nor2_0 U4 ( .x(n1), .a(bare_i), .b(force_bare) );
    aoi21_1 U6 ( .x(n2), .a(n3), .b(im_i), .c(r_h[1]) );
    inv_0 U8 ( .x(n3), .a(force_bare) );
    nor2i_0 U9 ( .x(n15), .a(wish_i), .b(force_bare) );
    nor2i_0 U10 ( .x(n14), .a(dm_i), .b(force_bare) );
    inv_0 U11 ( .x(e_h[1]), .a(n1) );
    buf_1 U15 ( .x(n6), .a(ah[31]) );
    buf_1 U16 ( .x(n7), .a(al[31]) );
    nand2_2 U17 ( .x(\e_l[2] ), .a(n2), .b(n1) );
    buf_1 U18 ( .x(r_h[1]), .a(n14) );
    inv_2 U19 ( .x(\e_h[0] ), .a(n2) );
    buf_3 U20 ( .x(\e_l[3] ), .a(\r_l[0] ) );
    buf_3 U21 ( .x(\e_l[0] ), .a(\r_l[2] ) );
    nand2i_2 U22 ( .x(e_l[1]), .a(n12), .b(n2) );
    buf_1 U23 ( .x(e_h[2]), .a(n15) );
    buf_1 U24 ( .x(r_l[3]), .a(n15) );
    buf_1 U25 ( .x(n12), .a(n15) );
endmodule


module chain_selement_ga_4 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_0 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[1] , \c[0] ;
    chain_selement_ga_4 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_5 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_1 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[1] , \c[0] ;
    chain_selement_ga_5 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_6 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_2 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[1] , \c[0] ;
    chain_selement_ga_6 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_7 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_3 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[1] , \c[0] ;
    chain_selement_ga_7 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_77 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_tx_iport ( o, rtxack, e_h, e_l, noa, r_h, r_l, rtxreq );
output [4:0] o;
input  [3:0] e_h;
input  [3:0] e_l;
input  [3:0] r_h;
input  [3:0] r_l;
input  noa, rtxreq;
output rtxack;
    wire \net52[0] , \net52[1] , \net55[0] , \net55[1] , \r3[2] , \r3[1] , 
        \r3[0] , \r0[2] , \r0[1] , \r0[0] , \r2[2] , \r2[1] , \r2[0] , 
        \last[0] , \last[1] , \last[2] , \last[3] , \last[4] , \r1[2] , 
        \r1[1] , \r1[0] , net6, eopsym, net9, net11, net16, net33, net60, 
        net40, net47, net50, \I8/nb , \I8/na , \I11/nc , \I11/nb , \I11/na , 
        \I7_0_/U25/U1/clr , \I7_0_/U25/U1/ob , \I7_1_/U25/U1/clr , 
        \I7_1_/U25/U1/ob ;
    assign o[3] = 1'b0;
    assign o[2] = 1'b0;
    route_symbol_0 I0 ( .o({\r3[2] , \r3[1] , \r3[0] }), .txack(net33), 
        .txack_last(\last[4] ), .e({e_h[3], e_l[3]}), .oa(net60), .r({r_h[3], 
        r_l[3]}), .txreq(rtxreq) );
    route_symbol_1 I1 ( .o({\r2[2] , \r2[1] , \r2[0] }), .txack(net40), 
        .txack_last(\last[3] ), .e({e_h[2], e_l[2]}), .oa(net60), .r({r_h[2], 
        r_l[2]}), .txreq(net33) );
    route_symbol_2 I2 ( .o({\r1[2] , \r1[1] , \r1[0] }), .txack(net47), 
        .txack_last(\last[2] ), .e({e_h[1], e_l[1]}), .oa(net60), .r({r_h[1], 
        r_l[1]}), .txreq(net40) );
    route_symbol_3 I3 ( .o({\r0[2] , \r0[1] , \r0[0] }), .txack(net50), 
        .txack_last(\last[1] ), .e({e_h[0], e_l[0]}), .oa(net60), .r({r_h[0], 
        r_l[0]}), .txreq(net47) );
    chain_selement_ga_77 I9 ( .Aa(\last[0] ), .Br(eopsym), .Ar(net50), .Ba(
        net60) );
    nor3_1 \I8/U27  ( .x(\I8/nb ), .a(o[4]), .b(o[3]), .c(o[2]) );
    nor2_1 \I8/U26  ( .x(\I8/na ), .a(o[1]), .b(o[0]) );
    nand2_2 \I8/U29  ( .x(net60), .a(\I8/nb ), .b(\I8/na ) );
    or2_1 \I13_0_/U12  ( .x(\net55[1] ), .a(\r1[0] ), .b(\r0[0] ) );
    or2_1 \I13_1_/U12  ( .x(\net55[0] ), .a(\r1[1] ), .b(\r0[1] ) );
    or2_1 \I14_0_/U12  ( .x(\net52[1] ), .a(\r3[0] ), .b(\r2[0] ) );
    or2_1 \I14_1_/U12  ( .x(\net52[0] ), .a(\r3[1] ), .b(\r2[1] ) );
    nand3_1 \I11/U31  ( .x(rtxack), .a(\I11/nc ), .b(\I11/nb ), .c(\I11/na )
         );
    inv_1 \I11/U33  ( .x(\I11/nc ), .a(\last[0] ) );
    nor2_1 \I11/U26  ( .x(\I11/na ), .a(\last[3] ), .b(\last[4] ) );
    nor2_1 \I11/U32  ( .x(\I11/nb ), .a(\last[1] ), .b(\last[2] ) );
    nor2_1 \I16/U5  ( .x(net16), .a(\r1[2] ), .b(\r0[2] ) );
    nor2_1 \I5/U5  ( .x(net11), .a(\r3[2] ), .b(\r2[2] ) );
    nand3_1 \I17/U9  ( .x(net9), .a(net6), .b(net11), .c(net16) );
    inv_1 \I18/U3  ( .x(net6), .a(eopsym) );
    oa31_1 \I7_0_/U25/U1/Uclr  ( .x(\I7_0_/U25/U1/clr ), .a(noa), .b(
        \net55[1] ), .c(\net52[1] ), .d(o[0]) );
    oaoi211_1 \I7_0_/U25/U1/Uaoi  ( .x(\I7_0_/U25/U1/ob ), .a(\net55[1] ), .b(
        \net52[1] ), .c(noa), .d(\I7_0_/U25/U1/clr ) );
    inv_2 \I7_0_/U25/U1/Ui  ( .x(o[0]), .a(\I7_0_/U25/U1/ob ) );
    oa31_1 \I7_1_/U25/U1/Uclr  ( .x(\I7_1_/U25/U1/clr ), .a(noa), .b(
        \net55[0] ), .c(\net52[0] ), .d(o[1]) );
    oaoi211_1 \I7_1_/U25/U1/Uaoi  ( .x(\I7_1_/U25/U1/ob ), .a(\net55[0] ), .b(
        \net52[0] ), .c(noa), .d(\I7_1_/U25/U1/clr ) );
    inv_2 \I7_1_/U25/U1/Ui  ( .x(o[1]), .a(\I7_1_/U25/U1/ob ) );
    ao222_1 \I15/U18/U1/U1  ( .x(o[4]), .a(noa), .b(net9), .c(noa), .d(o[4]), 
        .e(net9), .f(o[4]) );
endmodule


module chain_dr8bit_completion_16 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_17 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_18 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_19 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr32bit_completion_2 ( o, i );
input  [63:0] i;
output o;
    wire nx, \cd[3] , \cd[2] , ny, \cd[0] , \cd[1] , \U16/Z , \U6/Z , \U15/Z ;
    chain_dr8bit_completion_16 U11 ( .o(\cd[3] ), .i({i[63], i[62], i[61], 
        i[60], i[59], i[58], i[57], i[56], i[31], i[30], i[29], i[28], i[27], 
        i[26], i[25], i[24]}) );
    chain_dr8bit_completion_19 U14 ( .o(\cd[2] ), .i({i[55], i[54], i[53], 
        i[52], i[51], i[50], i[49], i[48], i[23], i[22], i[21], i[20], i[19], 
        i[18], i[17], i[16]}) );
    chain_dr8bit_completion_18 U13 ( .o(\cd[1] ), .i({i[47], i[46], i[45], 
        i[44], i[43], i[42], i[41], i[40], i[15], i[14], i[13], i[12], i[11], 
        i[10], i[9], i[8]}) );
    chain_dr8bit_completion_17 U12 ( .o(\cd[0] ), .i({i[39], i[38], i[37], 
        i[36], i[35], i[34], i[33], i[32], i[7], i[6], i[5], i[4], i[3], i[2], 
        i[1], i[0]}) );
    aoi222_1 \U16/U30/U1  ( .x(ny), .a(\cd[0] ), .b(\cd[1] ), .c(\cd[0] ), .d(
        \U16/Z ), .e(\cd[1] ), .f(\U16/Z ) );
    inv_1 \U16/U30/Uinv  ( .x(\U16/Z ), .a(ny) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(ny), .b(nx), .c(ny), .d(\U6/Z ), .e(nx), 
        .f(\U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U15/U30/U1  ( .x(nx), .a(\cd[3] ), .b(\cd[2] ), .c(\cd[3] ), .d(
        \U15/Z ), .e(\cd[2] ), .f(\U15/Z ) );
    inv_1 \U15/U30/Uinv  ( .x(\U15/Z ), .a(nx) );
endmodule


module chain_dr8bit_completion_20 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_21 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_22 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_23 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr32bit_completion_3 ( o, i );
input  [63:0] i;
output o;
    wire nx, \cd[3] , \cd[2] , ny, \cd[0] , \cd[1] , \U16/Z , \U6/Z , \U15/Z ;
    chain_dr8bit_completion_20 U11 ( .o(\cd[3] ), .i({i[63], i[62], i[61], 
        i[60], i[59], i[58], i[57], i[56], i[31], i[30], i[29], i[28], i[27], 
        i[26], i[25], i[24]}) );
    chain_dr8bit_completion_23 U14 ( .o(\cd[2] ), .i({i[55], i[54], i[53], 
        i[52], i[51], i[50], i[49], i[48], i[23], i[22], i[21], i[20], i[19], 
        i[18], i[17], i[16]}) );
    chain_dr8bit_completion_22 U13 ( .o(\cd[1] ), .i({i[47], i[46], i[45], 
        i[44], i[43], i[42], i[41], i[40], i[15], i[14], i[13], i[12], i[11], 
        i[10], i[9], i[8]}) );
    chain_dr8bit_completion_21 U12 ( .o(\cd[0] ), .i({i[39], i[38], i[37], 
        i[36], i[35], i[34], i[33], i[32], i[7], i[6], i[5], i[4], i[3], i[2], 
        i[1], i[0]}) );
    aoi222_1 \U16/U30/U1  ( .x(ny), .a(\cd[0] ), .b(\cd[1] ), .c(\cd[0] ), .d(
        \U16/Z ), .e(\cd[1] ), .f(\U16/Z ) );
    inv_1 \U16/U30/Uinv  ( .x(\U16/Z ), .a(ny) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(ny), .b(nx), .c(ny), .d(\U6/Z ), .e(nx), 
        .f(\U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U15/U30/U1  ( .x(nx), .a(\cd[3] ), .b(\cd[2] ), .c(\cd[3] ), .d(
        \U15/Z ), .e(\cd[2] ), .f(\U15/Z ) );
    inv_1 \U15/U30/Uinv  ( .x(\U15/Z ), .a(nx) );
endmodule


module chain_dr8bit_completion_50 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_51 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_selement_ga_32 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_33 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_34 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_35 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_36 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_37 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_38 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_39 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_40 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_41 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_icmux_0 ( ack, chainh, chainl, sendack, addr, col, itag, lock, 
    nReset, nia, pred, rnw, sendreq, seq, size, wd );
output [7:0] chainh;
output [7:0] chainl;
input  [63:0] addr;
input  [5:0] col;
input  [9:0] itag;
input  [1:0] lock;
input  [1:0] pred;
input  [1:0] rnw;
input  [1:0] seq;
input  [3:0] size;
input  [63:0] wd;
input  nReset, nia, sendreq;
output ack, sendack;
    wire \net207[0] , \net207[1] , \net207[2] , \net207[3] , \net207[4] , 
        \net207[5] , \net207[6] , \net207[7] , \net207[8] , \net207[9] , 
        \net207[10] , \net207[11] , \net207[12] , \net207[13] , \net207[14] , 
        \net207[15] , \bs[0] , \bs[1] , \bs[2] , \bs[3] , \bs[4] , \bs[5] , 
        \bs[6] , \bs[7] , \bs[8] , \net231[0] , \net231[1] , \net231[2] , 
        \net231[3] , \net231[4] , \net231[5] , \net231[6] , \net231[7] , 
        \net231[8] , \net231[9] , \net231[10] , \net231[11] , \net231[12] , 
        \net231[13] , \net231[14] , \net231[15] , \hdr[4] , \net234[0] , 
        \net234[1] , \net234[2] , \net234[3] , \net234[4] , \net234[5] , 
        \net234[6] , \net234[7] , \net234[8] , \net234[9] , \net234[10] , 
        \net234[11] , \net234[12] , \net234[13] , \net234[14] , \net234[15] , 
        \net217[0] , \net217[1] , \net217[2] , \net217[3] , \net217[4] , 
        \net217[5] , \net217[6] , \net217[7] , \net217[8] , \net217[9] , 
        \net217[10] , \net217[11] , \net217[12] , \net217[13] , \net217[14] , 
        \net217[15] , \net246[0] , \net246[1] , \net246[2] , \net246[3] , 
        \net246[4] , \net246[5] , \net246[6] , \net246[7] , \net246[8] , 
        \net246[9] , \net246[10] , \net246[11] , \net246[12] , \net246[13] , 
        \net246[14] , \net246[15] , \net243[0] , \net243[1] , \net243[2] , 
        \net243[3] , \net243[4] , \net243[5] , \net243[6] , \net243[7] , 
        \net243[8] , \net243[9] , \net243[10] , \net243[11] , \net243[12] , 
        \net243[13] , \net243[14] , \net243[15] , \net240[0] , \net240[1] , 
        \net240[2] , \net240[3] , \net240[4] , \net240[5] , \net240[6] , 
        \net240[7] , \net240[8] , \net240[9] , \net240[10] , \net240[11] , 
        \net240[12] , \net240[13] , \net240[14] , \net240[15] , \net219[0] , 
        \net219[1] , \net219[2] , \net219[3] , \net219[4] , \net219[5] , 
        \net219[6] , \net219[7] , \net219[8] , \net219[9] , \net219[10] , 
        \net219[11] , \net219[12] , \net219[13] , \net219[14] , \net219[15] , 
        \net237[0] , \net237[1] , \net237[2] , \net237[5] , \net237[6] , 
        \net237[7] , \net237[8] , \net237[9] , \net237[10] , \net237[11] , 
        \net237[12] , \net237[13] , \net237[14] , \net237[15] , \net222[0] , 
        \net222[1] , \net222[2] , \net222[3] , \net222[4] , \net222[5] , 
        \net222[6] , \net222[7] , \net222[8] , \net222[9] , \net222[10] , 
        \net222[11] , \net222[12] , \net222[13] , \net222[14] , \net222[15] , 
        \net225[0] , \net225[1] , \net225[2] , \net225[3] , \net225[4] , 
        \net225[5] , \net225[6] , \net225[7] , \net225[8] , \net225[9] , 
        \net225[10] , \net225[11] , \net225[12] , \net225[13] , \net225[14] , 
        \net225[15] , \net228[0] , \net228[1] , \net228[2] , \net228[3] , 
        \net228[4] , \net228[5] , \net228[6] , \net228[7] , \net228[8] , 
        \net228[9] , \net228[10] , \net228[11] , \net228[12] , \net228[13] , 
        \net228[14] , \net228[15] , \net212[0] , \net212[1] , \net212[2] , 
        \net212[3] , \net212[4] , \net212[5] , \net212[6] , \net212[7] , 
        \net212[8] , \net212[9] , \net212[10] , \net212[11] , \net212[12] , 
        \net212[13] , \net212[14] , \net212[15] , net138, net198, net176, 
        net132, net131, net136, net185, net187, net191, net293, net152, net146, 
        net148, net156, net160, net168, net172, net164, net289, net180, net189, 
        net249, net261, net251, net255, net253, net259, net269, net267, net263, 
        net265, \U40_0_/n5 , \U40_0_/n3 , \U40_0_/n4 , \U40_1_/n5 , 
        \U40_1_/n3 , \U40_1_/n4 , \U40_2_/n5 , \U40_2_/n3 , \U40_2_/n4 , 
        \U40_3_/n5 , \U40_3_/n3 , \U40_3_/n4 , \U40_4_/n5 , \U40_4_/n3 , 
        \U40_4_/n4 , \U40_5_/n5 , \U40_5_/n3 , \U40_5_/n4 , \U40_6_/n5 , 
        \U40_6_/n3 , \U40_6_/n4 , \U40_7_/n5 , \U40_7_/n3 , \U40_7_/n4 , 
        \U40_8_/n5 , \U40_8_/n3 , \U40_8_/n4 , \U40_9_/n5 , \U40_9_/n3 , 
        \U40_9_/n4 , \U40_10_/n5 , \U40_10_/n3 , \U40_10_/n4 , \U40_11_/n5 , 
        \U40_11_/n3 , \U40_11_/n4 , \U40_12_/n5 , \U40_12_/n3 , \U40_12_/n4 , 
        \U40_13_/n5 , \U40_13_/n3 , \U40_13_/n4 , \U40_14_/n5 , \U40_14_/n3 , 
        \U40_14_/n4 , \U40_15_/n5 , \U40_15_/n3 , \U40_15_/n4 , \U14_0_/n5 , 
        \U14_0_/n1 , \U14_0_/n2 , \U14_0_/n3 , \U14_0_/n4 , \U14_1_/n5 , 
        \U14_1_/n1 , \U14_1_/n2 , \U14_1_/n3 , \U14_1_/n4 , \U14_2_/n5 , 
        \U14_2_/n1 , \U14_2_/n2 , \U14_2_/n3 , \U14_2_/n4 , \U14_3_/n5 , 
        \U14_3_/n1 , \U14_3_/n2 , \U14_3_/n3 , \U14_3_/n4 , \U14_4_/n5 , 
        \U14_4_/n1 , \U14_4_/n2 , \U14_4_/n3 , \U14_4_/n4 , \U14_5_/n5 , 
        \U14_5_/n1 , \U14_5_/n2 , \U14_5_/n3 , \U14_5_/n4 , \U14_6_/n5 , 
        \U14_6_/n1 , \U14_6_/n2 , \U14_6_/n3 , \U14_6_/n4 , \U14_7_/n5 , 
        \U14_7_/n1 , \U14_7_/n2 , \U14_7_/n3 , \U14_7_/n4 , \U14_8_/n5 , 
        \U14_8_/n1 , \U14_8_/n2 , \U14_8_/n3 , \U14_8_/n4 , \U14_9_/n5 , 
        \U14_9_/n1 , \U14_9_/n2 , \U14_9_/n3 , \U14_9_/n4 , \U14_10_/n5 , 
        \U14_10_/n1 , \U14_10_/n2 , \U14_10_/n3 , \U14_10_/n4 , \U14_11_/n5 , 
        \U14_11_/n1 , \U14_11_/n2 , \U14_11_/n4 , \U14_12_/n5 , \U14_12_/n1 , 
        \U14_12_/n2 , \U14_12_/n4 , \U14_13_/n5 , \U14_13_/n1 , \U14_13_/n2 , 
        \U14_13_/n3 , \U14_13_/n4 , \U14_14_/n5 , \U14_14_/n1 , \U14_14_/n2 , 
        \U14_14_/n3 , \U14_14_/n4 , \U14_15_/n5 , \U14_15_/n1 , \U14_15_/n2 , 
        \U14_15_/n3 , \U14_15_/n4 , \U91_0_/n5 , \U91_0_/n1 , \U91_0_/n2 , 
        \U91_0_/n3 , \U91_0_/n4 , \U91_1_/n5 , \U91_1_/n1 , \U91_1_/n2 , 
        \U91_1_/n3 , \U91_1_/n4 , \U91_2_/n5 , \U91_2_/n1 , \U91_2_/n2 , 
        \U91_2_/n3 , \U91_2_/n4 , \U91_3_/n5 , \U91_3_/n1 , \U91_3_/n2 , 
        \U91_3_/n3 , \U91_3_/n4 , \U91_4_/n5 , \U91_4_/n1 , \U91_4_/n2 , 
        \U91_4_/n3 , \U91_4_/n4 , \U91_5_/n5 , \U91_5_/n1 , \U91_5_/n2 , 
        \U91_5_/n3 , \U91_5_/n4 , \U91_6_/n5 , \U91_6_/n1 , \U91_6_/n2 , 
        \U91_6_/n3 , \U91_6_/n4 , \U91_7_/n5 , \U91_7_/n1 , \U91_7_/n2 , 
        \U91_7_/n3 , \U91_7_/n4 , \U91_8_/n5 , \U91_8_/n1 , \U91_8_/n2 , 
        \U91_8_/n3 , \U91_8_/n4 , \U91_9_/n5 , \U91_9_/n1 , \U91_9_/n2 , 
        \U91_9_/n3 , \U91_9_/n4 , \U91_10_/n5 , \U91_10_/n1 , \U91_10_/n2 , 
        \U91_10_/n3 , \U91_10_/n4 , \U91_11_/n5 , \U91_11_/n1 , \U91_11_/n2 , 
        \U91_11_/n3 , \U91_11_/n4 , \U91_12_/n5 , \U91_12_/n1 , \U91_12_/n2 , 
        \U91_12_/n3 , \U91_12_/n4 , \U91_13_/n5 , \U91_13_/n1 , \U91_13_/n2 , 
        \U91_13_/n3 , \U91_13_/n4 , \U91_14_/n5 , \U91_14_/n1 , \U91_14_/n2 , 
        \U91_14_/n3 , \U91_14_/n4 , \U91_15_/n5 , \U91_15_/n1 , \U91_15_/n2 , 
        \U91_15_/n3 , \U91_15_/n4 , \U148/U21/nr , \U148/U21/nd , 
        \U148/U21/n2 , \U151/Z , n1;
    chain_selement_ga_33 U163 ( .Aa(net152), .Br(net146), .Ar(net148), .Ba(n1)
         );
    chain_selement_ga_34 U164 ( .Aa(net156), .Br(\bs[1] ), .Ar(net152), .Ba(
        net138) );
    chain_selement_ga_35 U165 ( .Aa(net160), .Br(\bs[2] ), .Ar(net156), .Ba(n1
        ) );
    chain_selement_ga_36 U166 ( .Aa(net168), .Br(\bs[3] ), .Ar(net160), .Ba(
        net138) );
    chain_selement_ga_40 U170 ( .Aa(net172), .Br(\bs[7] ), .Ar(net164), .Ba(
        net138) );
    chain_selement_ga_37 U167 ( .Aa(net132), .Br(\bs[4] ), .Ar(net168), .Ba(
        net138) );
    chain_selement_ga_41 U171 ( .Aa(net289), .Br(\bs[8] ), .Ar(net172), .Ba(
        net138) );
    chain_selement_ga_38 U168 ( .Aa(net180), .Br(\bs[5] ), .Ar(net176), .Ba(
        net138) );
    chain_selement_ga_39 U169 ( .Aa(net164), .Br(\bs[6] ), .Ar(net180), .Ba(n1
        ) );
    chain_selement_ga_32 U161 ( .Aa(net148), .Br(\bs[0] ), .Ar(\hdr[4] ), .Ba(
        n1) );
    chain_dr8bit_completion_50 U119 ( .o(net185), .i({col[5], col[4], col[3], 
        itag[9], itag[8], itag[7], itag[6], itag[5], col[2], col[1], col[0], 
        itag[4], itag[3], itag[2], itag[1], itag[0]}) );
    chain_dr8bit_completion_51 U147 ( .o(net187), .i({size[3], size[2], rnw[1], 
        1'b0, 1'b0, lock[1], pred[1], seq[1], size[1], size[0], rnw[0], 
        \hdr[4] , \hdr[4] , lock[0], pred[0], seq[0]}) );
    chain_dr32bit_completion_2 U117 ( .o(net189), .i(wd) );
    chain_dr32bit_completion_3 U118 ( .o(net191), .i(addr) );
    or2_4 \U122/U12  ( .x(net293), .a(net189), .b(net131) );
    or2_4 \U53/U12  ( .x(sendack), .a(net131), .b(net289) );
    and2_1 \U32_0_/U8  ( .x(\net246[15] ), .a(itag[0]), .b(net265) );
    and2_1 \U32_1_/U8  ( .x(\net246[14] ), .a(itag[1]), .b(net265) );
    and2_1 \U32_2_/U8  ( .x(\net246[13] ), .a(itag[2]), .b(net265) );
    and2_1 \U32_3_/U8  ( .x(\net246[12] ), .a(itag[3]), .b(net265) );
    and2_1 \U32_4_/U8  ( .x(\net246[11] ), .a(itag[4]), .b(net265) );
    and2_1 \U32_5_/U8  ( .x(\net246[10] ), .a(col[0]), .b(net265) );
    and2_1 \U32_6_/U8  ( .x(\net246[9] ), .a(col[1]), .b(net265) );
    and2_1 \U32_7_/U8  ( .x(\net246[8] ), .a(col[2]), .b(net265) );
    and2_1 \U32_8_/U8  ( .x(\net246[7] ), .a(itag[5]), .b(net265) );
    and2_1 \U32_9_/U8  ( .x(\net246[6] ), .a(itag[6]), .b(net265) );
    and2_1 \U32_10_/U8  ( .x(\net246[5] ), .a(itag[7]), .b(net265) );
    and2_1 \U32_11_/U8  ( .x(\net246[4] ), .a(itag[8]), .b(net265) );
    and2_1 \U32_12_/U8  ( .x(\net246[3] ), .a(itag[9]), .b(net265) );
    and2_1 \U32_13_/U8  ( .x(\net246[2] ), .a(col[3]), .b(net265) );
    and2_1 \U32_14_/U8  ( .x(\net246[1] ), .a(col[4]), .b(net265) );
    and2_1 \U32_15_/U8  ( .x(\net246[0] ), .a(col[5]), .b(net265) );
    and2_1 \U76_0_/U8  ( .x(\net243[15] ), .a(wd[8]), .b(net263) );
    and2_1 \U76_1_/U8  ( .x(\net243[14] ), .a(wd[9]), .b(net263) );
    and2_1 \U76_2_/U8  ( .x(\net243[13] ), .a(wd[10]), .b(net263) );
    and2_1 \U76_3_/U8  ( .x(\net243[12] ), .a(wd[11]), .b(net263) );
    and2_1 \U76_4_/U8  ( .x(\net243[11] ), .a(wd[12]), .b(net263) );
    and2_1 \U76_5_/U8  ( .x(\net243[10] ), .a(wd[13]), .b(net263) );
    and2_1 \U76_6_/U8  ( .x(\net243[9] ), .a(wd[14]), .b(net263) );
    and2_1 \U76_7_/U8  ( .x(\net243[8] ), .a(wd[15]), .b(net263) );
    and2_1 \U76_8_/U8  ( .x(\net243[7] ), .a(wd[40]), .b(net263) );
    and2_1 \U76_9_/U8  ( .x(\net243[6] ), .a(wd[41]), .b(net263) );
    and2_1 \U76_10_/U8  ( .x(\net243[5] ), .a(wd[42]), .b(net263) );
    and2_1 \U76_11_/U8  ( .x(\net243[4] ), .a(wd[43]), .b(net263) );
    and2_1 \U76_12_/U8  ( .x(\net243[3] ), .a(wd[44]), .b(net263) );
    and2_1 \U76_13_/U8  ( .x(\net243[2] ), .a(wd[45]), .b(net263) );
    and2_1 \U76_14_/U8  ( .x(\net243[1] ), .a(wd[46]), .b(net263) );
    and2_1 \U76_15_/U8  ( .x(\net243[0] ), .a(wd[47]), .b(net263) );
    and2_1 \U80_0_/U8  ( .x(\net240[15] ), .a(wd[16]), .b(net267) );
    and2_1 \U80_1_/U8  ( .x(\net240[14] ), .a(wd[17]), .b(net267) );
    and2_1 \U80_2_/U8  ( .x(\net240[13] ), .a(wd[18]), .b(net267) );
    and2_1 \U80_3_/U8  ( .x(\net240[12] ), .a(wd[19]), .b(net267) );
    and2_1 \U80_4_/U8  ( .x(\net240[11] ), .a(wd[20]), .b(net267) );
    and2_1 \U80_5_/U8  ( .x(\net240[10] ), .a(wd[21]), .b(net267) );
    and2_1 \U80_6_/U8  ( .x(\net240[9] ), .a(wd[22]), .b(net267) );
    and2_1 \U80_7_/U8  ( .x(\net240[8] ), .a(wd[23]), .b(net267) );
    and2_1 \U80_8_/U8  ( .x(\net240[7] ), .a(wd[48]), .b(net267) );
    and2_1 \U80_9_/U8  ( .x(\net240[6] ), .a(wd[49]), .b(net267) );
    and2_1 \U80_10_/U8  ( .x(\net240[5] ), .a(wd[50]), .b(net267) );
    and2_1 \U80_11_/U8  ( .x(\net240[4] ), .a(wd[51]), .b(net267) );
    and2_1 \U80_12_/U8  ( .x(\net240[3] ), .a(wd[52]), .b(net267) );
    and2_1 \U80_13_/U8  ( .x(\net240[2] ), .a(wd[53]), .b(net267) );
    and2_1 \U80_14_/U8  ( .x(\net240[1] ), .a(wd[54]), .b(net267) );
    and2_1 \U80_15_/U8  ( .x(\net240[0] ), .a(wd[55]), .b(net267) );
    and2_1 \U128_0_/U8  ( .x(\net237[15] ), .a(seq[0]), .b(net269) );
    and2_1 \U128_1_/U8  ( .x(\net237[14] ), .a(pred[0]), .b(net269) );
    and2_1 \U128_2_/U8  ( .x(\net237[13] ), .a(lock[0]), .b(net269) );
    and2_1 \U128_3_/U8  ( .x(\net237[12] ), .a(\hdr[4] ), .b(net269) );
    and2_1 \U128_4_/U8  ( .x(\net237[11] ), .a(\hdr[4] ), .b(net269) );
    and2_1 \U128_5_/U8  ( .x(\net237[10] ), .a(rnw[0]), .b(net269) );
    and2_1 \U128_6_/U8  ( .x(\net237[9] ), .a(size[0]), .b(net269) );
    and2_1 \U128_7_/U8  ( .x(\net237[8] ), .a(size[1]), .b(net269) );
    and2_1 \U128_8_/U8  ( .x(\net237[7] ), .a(seq[1]), .b(net269) );
    and2_1 \U128_9_/U8  ( .x(\net237[6] ), .a(pred[1]), .b(net269) );
    and2_1 \U128_10_/U8  ( .x(\net237[5] ), .a(lock[1]), .b(net269) );
    and2_1 \U128_13_/U8  ( .x(\net237[2] ), .a(rnw[1]), .b(net269) );
    and2_1 \U128_14_/U8  ( .x(\net237[1] ), .a(size[2]), .b(net269) );
    and2_1 \U128_15_/U8  ( .x(\net237[0] ), .a(size[3]), .b(net269) );
    and2_1 \U37_0_/U8  ( .x(\net234[15] ), .a(addr[8]), .b(net259) );
    and2_1 \U37_1_/U8  ( .x(\net234[14] ), .a(addr[9]), .b(net259) );
    and2_1 \U37_2_/U8  ( .x(\net234[13] ), .a(addr[10]), .b(net259) );
    and2_1 \U37_3_/U8  ( .x(\net234[12] ), .a(addr[11]), .b(net259) );
    and2_1 \U37_4_/U8  ( .x(\net234[11] ), .a(addr[12]), .b(net259) );
    and2_1 \U37_5_/U8  ( .x(\net234[10] ), .a(addr[13]), .b(net259) );
    and2_1 \U37_6_/U8  ( .x(\net234[9] ), .a(addr[14]), .b(net259) );
    and2_1 \U37_7_/U8  ( .x(\net234[8] ), .a(addr[15]), .b(net259) );
    and2_1 \U37_8_/U8  ( .x(\net234[7] ), .a(addr[40]), .b(net259) );
    and2_1 \U37_9_/U8  ( .x(\net234[6] ), .a(addr[41]), .b(net259) );
    and2_1 \U37_10_/U8  ( .x(\net234[5] ), .a(addr[42]), .b(net259) );
    and2_1 \U37_11_/U8  ( .x(\net234[4] ), .a(addr[43]), .b(net259) );
    and2_1 \U37_12_/U8  ( .x(\net234[3] ), .a(addr[44]), .b(net259) );
    and2_1 \U37_13_/U8  ( .x(\net234[2] ), .a(addr[45]), .b(net259) );
    and2_1 \U37_14_/U8  ( .x(\net234[1] ), .a(addr[46]), .b(net259) );
    and2_1 \U37_15_/U8  ( .x(\net234[0] ), .a(addr[47]), .b(net259) );
    and2_1 \U33_0_/U8  ( .x(\net231[15] ), .a(addr[16]), .b(net253) );
    and2_1 \U33_1_/U8  ( .x(\net231[14] ), .a(addr[17]), .b(net253) );
    and2_1 \U33_2_/U8  ( .x(\net231[13] ), .a(addr[18]), .b(net253) );
    and2_1 \U33_3_/U8  ( .x(\net231[12] ), .a(addr[19]), .b(net253) );
    and2_1 \U33_4_/U8  ( .x(\net231[11] ), .a(addr[20]), .b(net253) );
    and2_1 \U33_5_/U8  ( .x(\net231[10] ), .a(addr[21]), .b(net253) );
    and2_1 \U33_6_/U8  ( .x(\net231[9] ), .a(addr[22]), .b(net253) );
    and2_1 \U33_7_/U8  ( .x(\net231[8] ), .a(addr[23]), .b(net253) );
    and2_1 \U33_8_/U8  ( .x(\net231[7] ), .a(addr[48]), .b(net253) );
    and2_1 \U33_9_/U8  ( .x(\net231[6] ), .a(addr[49]), .b(net253) );
    and2_1 \U33_10_/U8  ( .x(\net231[5] ), .a(addr[50]), .b(net253) );
    and2_1 \U33_11_/U8  ( .x(\net231[4] ), .a(addr[51]), .b(net253) );
    and2_1 \U33_12_/U8  ( .x(\net231[3] ), .a(addr[52]), .b(net253) );
    and2_1 \U33_13_/U8  ( .x(\net231[2] ), .a(addr[53]), .b(net253) );
    and2_1 \U33_14_/U8  ( .x(\net231[1] ), .a(addr[54]), .b(net253) );
    and2_1 \U33_15_/U8  ( .x(\net231[0] ), .a(addr[55]), .b(net253) );
    and2_1 \U81_0_/U8  ( .x(\net228[15] ), .a(wd[24]), .b(net255) );
    and2_1 \U81_1_/U8  ( .x(\net228[14] ), .a(wd[25]), .b(net255) );
    and2_1 \U81_2_/U8  ( .x(\net228[13] ), .a(wd[26]), .b(net255) );
    and2_1 \U81_3_/U8  ( .x(\net228[12] ), .a(wd[27]), .b(net255) );
    and2_1 \U81_4_/U8  ( .x(\net228[11] ), .a(wd[28]), .b(net255) );
    and2_1 \U81_5_/U8  ( .x(\net228[10] ), .a(wd[29]), .b(net255) );
    and2_1 \U81_6_/U8  ( .x(\net228[9] ), .a(wd[30]), .b(net255) );
    and2_1 \U81_7_/U8  ( .x(\net228[8] ), .a(wd[31]), .b(net255) );
    and2_1 \U81_8_/U8  ( .x(\net228[7] ), .a(wd[56]), .b(net255) );
    and2_1 \U81_9_/U8  ( .x(\net228[6] ), .a(wd[57]), .b(net255) );
    and2_1 \U81_10_/U8  ( .x(\net228[5] ), .a(wd[58]), .b(net255) );
    and2_1 \U81_11_/U8  ( .x(\net228[4] ), .a(wd[59]), .b(net255) );
    and2_1 \U81_12_/U8  ( .x(\net228[3] ), .a(wd[60]), .b(net255) );
    and2_1 \U81_13_/U8  ( .x(\net228[2] ), .a(wd[61]), .b(net255) );
    and2_1 \U81_14_/U8  ( .x(\net228[1] ), .a(wd[62]), .b(net255) );
    and2_1 \U81_15_/U8  ( .x(\net228[0] ), .a(wd[63]), .b(net255) );
    and2_1 \U34_0_/U8  ( .x(\net225[15] ), .a(addr[0]), .b(net251) );
    and2_1 \U34_1_/U8  ( .x(\net225[14] ), .a(addr[1]), .b(net251) );
    and2_1 \U34_2_/U8  ( .x(\net225[13] ), .a(addr[2]), .b(net251) );
    and2_1 \U34_3_/U8  ( .x(\net225[12] ), .a(addr[3]), .b(net251) );
    and2_1 \U34_4_/U8  ( .x(\net225[11] ), .a(addr[4]), .b(net251) );
    and2_1 \U34_5_/U8  ( .x(\net225[10] ), .a(addr[5]), .b(net251) );
    and2_1 \U34_6_/U8  ( .x(\net225[9] ), .a(addr[6]), .b(net251) );
    and2_1 \U34_7_/U8  ( .x(\net225[8] ), .a(addr[7]), .b(net251) );
    and2_1 \U34_8_/U8  ( .x(\net225[7] ), .a(addr[32]), .b(net251) );
    and2_1 \U34_9_/U8  ( .x(\net225[6] ), .a(addr[33]), .b(net251) );
    and2_1 \U34_10_/U8  ( .x(\net225[5] ), .a(addr[34]), .b(net251) );
    and2_1 \U34_11_/U8  ( .x(\net225[4] ), .a(addr[35]), .b(net251) );
    and2_1 \U34_12_/U8  ( .x(\net225[3] ), .a(addr[36]), .b(net251) );
    and2_1 \U34_13_/U8  ( .x(\net225[2] ), .a(addr[37]), .b(net251) );
    and2_1 \U34_14_/U8  ( .x(\net225[1] ), .a(addr[38]), .b(net251) );
    and2_1 \U34_15_/U8  ( .x(\net225[0] ), .a(addr[39]), .b(net251) );
    and2_1 \U30_0_/U8  ( .x(\net222[15] ), .a(addr[24]), .b(net261) );
    and2_1 \U30_1_/U8  ( .x(\net222[14] ), .a(addr[25]), .b(net261) );
    and2_1 \U30_2_/U8  ( .x(\net222[13] ), .a(addr[26]), .b(net261) );
    and2_1 \U30_3_/U8  ( .x(\net222[12] ), .a(addr[27]), .b(net261) );
    and2_1 \U30_4_/U8  ( .x(\net222[11] ), .a(addr[28]), .b(net261) );
    and2_1 \U30_5_/U8  ( .x(\net222[10] ), .a(addr[29]), .b(net261) );
    and2_1 \U30_6_/U8  ( .x(\net222[9] ), .a(addr[30]), .b(net261) );
    and2_1 \U30_7_/U8  ( .x(\net222[8] ), .a(addr[31]), .b(net261) );
    and2_1 \U30_8_/U8  ( .x(\net222[7] ), .a(addr[56]), .b(net261) );
    and2_1 \U30_9_/U8  ( .x(\net222[6] ), .a(addr[57]), .b(net261) );
    and2_1 \U30_10_/U8  ( .x(\net222[5] ), .a(addr[58]), .b(net261) );
    and2_1 \U30_11_/U8  ( .x(\net222[4] ), .a(addr[59]), .b(net261) );
    and2_1 \U30_12_/U8  ( .x(\net222[3] ), .a(addr[60]), .b(net261) );
    and2_1 \U30_13_/U8  ( .x(\net222[2] ), .a(addr[61]), .b(net261) );
    and2_1 \U30_14_/U8  ( .x(\net222[1] ), .a(addr[62]), .b(net261) );
    and2_1 \U30_15_/U8  ( .x(\net222[0] ), .a(addr[63]), .b(net261) );
    and2_1 \U82_0_/U8  ( .x(\net219[15] ), .a(wd[0]), .b(net249) );
    and2_1 \U82_1_/U8  ( .x(\net219[14] ), .a(wd[1]), .b(net249) );
    and2_1 \U82_2_/U8  ( .x(\net219[13] ), .a(wd[2]), .b(net249) );
    and2_1 \U82_3_/U8  ( .x(\net219[12] ), .a(wd[3]), .b(net249) );
    and2_1 \U82_4_/U8  ( .x(\net219[11] ), .a(wd[4]), .b(net249) );
    and2_1 \U82_5_/U8  ( .x(\net219[10] ), .a(wd[5]), .b(net249) );
    and2_1 \U82_6_/U8  ( .x(\net219[9] ), .a(wd[6]), .b(net249) );
    and2_1 \U82_7_/U8  ( .x(\net219[8] ), .a(wd[7]), .b(net249) );
    and2_1 \U82_8_/U8  ( .x(\net219[7] ), .a(wd[32]), .b(net249) );
    and2_1 \U82_9_/U8  ( .x(\net219[6] ), .a(wd[33]), .b(net249) );
    and2_1 \U82_10_/U8  ( .x(\net219[5] ), .a(wd[34]), .b(net249) );
    and2_1 \U82_11_/U8  ( .x(\net219[4] ), .a(wd[35]), .b(net249) );
    and2_1 \U82_12_/U8  ( .x(\net219[3] ), .a(wd[36]), .b(net249) );
    and2_1 \U82_13_/U8  ( .x(\net219[2] ), .a(wd[37]), .b(net249) );
    and2_1 \U82_14_/U8  ( .x(\net219[1] ), .a(wd[38]), .b(net249) );
    and2_1 \U82_15_/U8  ( .x(\net219[0] ), .a(wd[39]), .b(net249) );
    inv_1 \U40_0_/U3  ( .x(\U40_0_/n3 ), .a(\net225[15] ) );
    inv_1 \U40_0_/U4  ( .x(\U40_0_/n4 ), .a(\net234[15] ) );
    inv_1 \U40_0_/U5  ( .x(\net217[15] ), .a(\U40_0_/n5 ) );
    inv_1 \U40_1_/U3  ( .x(\U40_1_/n3 ), .a(\net225[14] ) );
    inv_1 \U40_1_/U4  ( .x(\U40_1_/n4 ), .a(\net234[14] ) );
    inv_1 \U40_1_/U5  ( .x(\net217[14] ), .a(\U40_1_/n5 ) );
    inv_1 \U40_2_/U3  ( .x(\U40_2_/n3 ), .a(\net225[13] ) );
    inv_1 \U40_2_/U4  ( .x(\U40_2_/n4 ), .a(\net234[13] ) );
    inv_1 \U40_2_/U5  ( .x(\net217[13] ), .a(\U40_2_/n5 ) );
    inv_1 \U40_3_/U3  ( .x(\U40_3_/n3 ), .a(\net225[12] ) );
    inv_1 \U40_3_/U4  ( .x(\U40_3_/n4 ), .a(\net234[12] ) );
    inv_1 \U40_3_/U5  ( .x(\net217[12] ), .a(\U40_3_/n5 ) );
    inv_1 \U40_4_/U3  ( .x(\U40_4_/n3 ), .a(\net225[11] ) );
    inv_1 \U40_4_/U4  ( .x(\U40_4_/n4 ), .a(\net234[11] ) );
    inv_1 \U40_4_/U5  ( .x(\net217[11] ), .a(\U40_4_/n5 ) );
    inv_1 \U40_5_/U3  ( .x(\U40_5_/n3 ), .a(\net225[10] ) );
    inv_1 \U40_5_/U4  ( .x(\U40_5_/n4 ), .a(\net234[10] ) );
    inv_1 \U40_5_/U5  ( .x(\net217[10] ), .a(\U40_5_/n5 ) );
    inv_1 \U40_6_/U3  ( .x(\U40_6_/n3 ), .a(\net225[9] ) );
    inv_1 \U40_6_/U4  ( .x(\U40_6_/n4 ), .a(\net234[9] ) );
    inv_1 \U40_6_/U5  ( .x(\net217[9] ), .a(\U40_6_/n5 ) );
    inv_1 \U40_7_/U3  ( .x(\U40_7_/n3 ), .a(\net225[8] ) );
    inv_1 \U40_7_/U4  ( .x(\U40_7_/n4 ), .a(\net234[8] ) );
    inv_1 \U40_7_/U5  ( .x(\net217[8] ), .a(\U40_7_/n5 ) );
    inv_1 \U40_8_/U3  ( .x(\U40_8_/n3 ), .a(\net225[7] ) );
    inv_1 \U40_8_/U4  ( .x(\U40_8_/n4 ), .a(\net234[7] ) );
    inv_1 \U40_8_/U5  ( .x(\net217[7] ), .a(\U40_8_/n5 ) );
    inv_1 \U40_9_/U3  ( .x(\U40_9_/n3 ), .a(\net225[6] ) );
    inv_1 \U40_9_/U4  ( .x(\U40_9_/n4 ), .a(\net234[6] ) );
    inv_1 \U40_9_/U5  ( .x(\net217[6] ), .a(\U40_9_/n5 ) );
    inv_1 \U40_10_/U3  ( .x(\U40_10_/n3 ), .a(\net225[5] ) );
    inv_1 \U40_10_/U4  ( .x(\U40_10_/n4 ), .a(\net234[5] ) );
    inv_1 \U40_10_/U5  ( .x(\net217[5] ), .a(\U40_10_/n5 ) );
    inv_1 \U40_11_/U3  ( .x(\U40_11_/n3 ), .a(\net225[4] ) );
    inv_1 \U40_11_/U4  ( .x(\U40_11_/n4 ), .a(\net234[4] ) );
    inv_1 \U40_11_/U5  ( .x(\net217[4] ), .a(\U40_11_/n5 ) );
    inv_1 \U40_12_/U3  ( .x(\U40_12_/n3 ), .a(\net225[3] ) );
    inv_1 \U40_12_/U4  ( .x(\U40_12_/n4 ), .a(\net234[3] ) );
    inv_1 \U40_12_/U5  ( .x(\net217[3] ), .a(\U40_12_/n5 ) );
    inv_1 \U40_13_/U3  ( .x(\U40_13_/n3 ), .a(\net225[2] ) );
    inv_1 \U40_13_/U4  ( .x(\U40_13_/n4 ), .a(\net234[2] ) );
    inv_1 \U40_13_/U5  ( .x(\net217[2] ), .a(\U40_13_/n5 ) );
    inv_1 \U40_14_/U3  ( .x(\U40_14_/n3 ), .a(\net225[1] ) );
    inv_1 \U40_14_/U4  ( .x(\U40_14_/n4 ), .a(\net234[1] ) );
    inv_1 \U40_14_/U5  ( .x(\net217[1] ), .a(\U40_14_/n5 ) );
    inv_1 \U40_15_/U3  ( .x(\U40_15_/n3 ), .a(\net225[0] ) );
    inv_1 \U40_15_/U4  ( .x(\U40_15_/n4 ), .a(\net234[0] ) );
    inv_1 \U40_15_/U5  ( .x(\net217[0] ), .a(\U40_15_/n5 ) );
    and4_1 \U14_0_/U16  ( .x(\U14_0_/n5 ), .a(\U14_0_/n1 ), .b(\U14_0_/n2 ), 
        .c(\U14_0_/n3 ), .d(\U14_0_/n4 ) );
    inv_1 \U14_0_/U1  ( .x(\U14_0_/n1 ), .a(\net231[15] ) );
    inv_1 \U14_0_/U2  ( .x(\U14_0_/n2 ), .a(\net222[15] ) );
    inv_1 \U14_0_/U3  ( .x(\U14_0_/n3 ), .a(\net237[15] ) );
    inv_1 \U14_0_/U4  ( .x(\U14_0_/n4 ), .a(\net246[15] ) );
    inv_1 \U14_0_/U5  ( .x(\net212[15] ), .a(\U14_0_/n5 ) );
    and4_1 \U14_1_/U16  ( .x(\U14_1_/n5 ), .a(\U14_1_/n1 ), .b(\U14_1_/n2 ), 
        .c(\U14_1_/n3 ), .d(\U14_1_/n4 ) );
    inv_1 \U14_1_/U1  ( .x(\U14_1_/n1 ), .a(\net231[14] ) );
    inv_1 \U14_1_/U2  ( .x(\U14_1_/n2 ), .a(\net222[14] ) );
    inv_1 \U14_1_/U3  ( .x(\U14_1_/n3 ), .a(\net237[14] ) );
    inv_1 \U14_1_/U4  ( .x(\U14_1_/n4 ), .a(\net246[14] ) );
    inv_1 \U14_1_/U5  ( .x(\net212[14] ), .a(\U14_1_/n5 ) );
    and4_1 \U14_2_/U16  ( .x(\U14_2_/n5 ), .a(\U14_2_/n1 ), .b(\U14_2_/n2 ), 
        .c(\U14_2_/n3 ), .d(\U14_2_/n4 ) );
    inv_1 \U14_2_/U1  ( .x(\U14_2_/n1 ), .a(\net231[13] ) );
    inv_1 \U14_2_/U2  ( .x(\U14_2_/n2 ), .a(\net222[13] ) );
    inv_1 \U14_2_/U3  ( .x(\U14_2_/n3 ), .a(\net237[13] ) );
    inv_1 \U14_2_/U4  ( .x(\U14_2_/n4 ), .a(\net246[13] ) );
    inv_1 \U14_2_/U5  ( .x(\net212[13] ), .a(\U14_2_/n5 ) );
    and4_1 \U14_3_/U16  ( .x(\U14_3_/n5 ), .a(\U14_3_/n1 ), .b(\U14_3_/n2 ), 
        .c(\U14_3_/n3 ), .d(\U14_3_/n4 ) );
    inv_1 \U14_3_/U1  ( .x(\U14_3_/n1 ), .a(\net231[12] ) );
    inv_1 \U14_3_/U2  ( .x(\U14_3_/n2 ), .a(\net222[12] ) );
    inv_1 \U14_3_/U3  ( .x(\U14_3_/n3 ), .a(\net237[12] ) );
    inv_1 \U14_3_/U4  ( .x(\U14_3_/n4 ), .a(\net246[12] ) );
    inv_1 \U14_3_/U5  ( .x(\net212[12] ), .a(\U14_3_/n5 ) );
    and4_1 \U14_4_/U16  ( .x(\U14_4_/n5 ), .a(\U14_4_/n1 ), .b(\U14_4_/n2 ), 
        .c(\U14_4_/n3 ), .d(\U14_4_/n4 ) );
    inv_1 \U14_4_/U1  ( .x(\U14_4_/n1 ), .a(\net231[11] ) );
    inv_1 \U14_4_/U2  ( .x(\U14_4_/n2 ), .a(\net222[11] ) );
    inv_1 \U14_4_/U3  ( .x(\U14_4_/n3 ), .a(\net237[11] ) );
    inv_1 \U14_4_/U4  ( .x(\U14_4_/n4 ), .a(\net246[11] ) );
    inv_1 \U14_4_/U5  ( .x(\net212[11] ), .a(\U14_4_/n5 ) );
    and4_1 \U14_5_/U16  ( .x(\U14_5_/n5 ), .a(\U14_5_/n1 ), .b(\U14_5_/n2 ), 
        .c(\U14_5_/n3 ), .d(\U14_5_/n4 ) );
    inv_1 \U14_5_/U1  ( .x(\U14_5_/n1 ), .a(\net231[10] ) );
    inv_1 \U14_5_/U2  ( .x(\U14_5_/n2 ), .a(\net222[10] ) );
    inv_1 \U14_5_/U3  ( .x(\U14_5_/n3 ), .a(\net237[10] ) );
    inv_1 \U14_5_/U4  ( .x(\U14_5_/n4 ), .a(\net246[10] ) );
    inv_1 \U14_5_/U5  ( .x(\net212[10] ), .a(\U14_5_/n5 ) );
    and4_1 \U14_6_/U16  ( .x(\U14_6_/n5 ), .a(\U14_6_/n1 ), .b(\U14_6_/n2 ), 
        .c(\U14_6_/n3 ), .d(\U14_6_/n4 ) );
    inv_1 \U14_6_/U1  ( .x(\U14_6_/n1 ), .a(\net231[9] ) );
    inv_1 \U14_6_/U2  ( .x(\U14_6_/n2 ), .a(\net222[9] ) );
    inv_1 \U14_6_/U3  ( .x(\U14_6_/n3 ), .a(\net237[9] ) );
    inv_1 \U14_6_/U4  ( .x(\U14_6_/n4 ), .a(\net246[9] ) );
    inv_1 \U14_6_/U5  ( .x(\net212[9] ), .a(\U14_6_/n5 ) );
    and4_1 \U14_7_/U16  ( .x(\U14_7_/n5 ), .a(\U14_7_/n1 ), .b(\U14_7_/n2 ), 
        .c(\U14_7_/n3 ), .d(\U14_7_/n4 ) );
    inv_1 \U14_7_/U1  ( .x(\U14_7_/n1 ), .a(\net231[8] ) );
    inv_1 \U14_7_/U2  ( .x(\U14_7_/n2 ), .a(\net222[8] ) );
    inv_1 \U14_7_/U3  ( .x(\U14_7_/n3 ), .a(\net237[8] ) );
    inv_1 \U14_7_/U4  ( .x(\U14_7_/n4 ), .a(\net246[8] ) );
    inv_1 \U14_7_/U5  ( .x(\net212[8] ), .a(\U14_7_/n5 ) );
    and4_1 \U14_8_/U16  ( .x(\U14_8_/n5 ), .a(\U14_8_/n1 ), .b(\U14_8_/n2 ), 
        .c(\U14_8_/n3 ), .d(\U14_8_/n4 ) );
    inv_1 \U14_8_/U1  ( .x(\U14_8_/n1 ), .a(\net231[7] ) );
    inv_1 \U14_8_/U2  ( .x(\U14_8_/n2 ), .a(\net222[7] ) );
    inv_1 \U14_8_/U3  ( .x(\U14_8_/n3 ), .a(\net237[7] ) );
    inv_1 \U14_8_/U4  ( .x(\U14_8_/n4 ), .a(\net246[7] ) );
    inv_1 \U14_8_/U5  ( .x(\net212[7] ), .a(\U14_8_/n5 ) );
    and4_1 \U14_9_/U16  ( .x(\U14_9_/n5 ), .a(\U14_9_/n1 ), .b(\U14_9_/n2 ), 
        .c(\U14_9_/n3 ), .d(\U14_9_/n4 ) );
    inv_1 \U14_9_/U1  ( .x(\U14_9_/n1 ), .a(\net231[6] ) );
    inv_1 \U14_9_/U2  ( .x(\U14_9_/n2 ), .a(\net222[6] ) );
    inv_1 \U14_9_/U3  ( .x(\U14_9_/n3 ), .a(\net237[6] ) );
    inv_1 \U14_9_/U4  ( .x(\U14_9_/n4 ), .a(\net246[6] ) );
    inv_1 \U14_9_/U5  ( .x(\net212[6] ), .a(\U14_9_/n5 ) );
    and4_1 \U14_10_/U16  ( .x(\U14_10_/n5 ), .a(\U14_10_/n1 ), .b(\U14_10_/n2 
        ), .c(\U14_10_/n3 ), .d(\U14_10_/n4 ) );
    inv_1 \U14_10_/U1  ( .x(\U14_10_/n1 ), .a(\net231[5] ) );
    inv_1 \U14_10_/U2  ( .x(\U14_10_/n2 ), .a(\net222[5] ) );
    inv_1 \U14_10_/U3  ( .x(\U14_10_/n3 ), .a(\net237[5] ) );
    inv_1 \U14_10_/U4  ( .x(\U14_10_/n4 ), .a(\net246[5] ) );
    inv_1 \U14_10_/U5  ( .x(\net212[5] ), .a(\U14_10_/n5 ) );
    inv_1 \U14_11_/U1  ( .x(\U14_11_/n1 ), .a(\net231[4] ) );
    inv_1 \U14_11_/U2  ( .x(\U14_11_/n2 ), .a(\net222[4] ) );
    inv_1 \U14_11_/U4  ( .x(\U14_11_/n4 ), .a(\net246[4] ) );
    inv_1 \U14_11_/U5  ( .x(\net212[4] ), .a(\U14_11_/n5 ) );
    inv_1 \U14_12_/U1  ( .x(\U14_12_/n1 ), .a(\net231[3] ) );
    inv_1 \U14_12_/U2  ( .x(\U14_12_/n2 ), .a(\net222[3] ) );
    inv_1 \U14_12_/U4  ( .x(\U14_12_/n4 ), .a(\net246[3] ) );
    inv_1 \U14_12_/U5  ( .x(\net212[3] ), .a(\U14_12_/n5 ) );
    and4_1 \U14_13_/U16  ( .x(\U14_13_/n5 ), .a(\U14_13_/n1 ), .b(\U14_13_/n2 
        ), .c(\U14_13_/n3 ), .d(\U14_13_/n4 ) );
    inv_1 \U14_13_/U1  ( .x(\U14_13_/n1 ), .a(\net231[2] ) );
    inv_1 \U14_13_/U2  ( .x(\U14_13_/n2 ), .a(\net222[2] ) );
    inv_1 \U14_13_/U3  ( .x(\U14_13_/n3 ), .a(\net237[2] ) );
    inv_1 \U14_13_/U4  ( .x(\U14_13_/n4 ), .a(\net246[2] ) );
    inv_1 \U14_13_/U5  ( .x(\net212[2] ), .a(\U14_13_/n5 ) );
    and4_1 \U14_14_/U16  ( .x(\U14_14_/n5 ), .a(\U14_14_/n1 ), .b(\U14_14_/n2 
        ), .c(\U14_14_/n3 ), .d(\U14_14_/n4 ) );
    inv_1 \U14_14_/U1  ( .x(\U14_14_/n1 ), .a(\net231[1] ) );
    inv_1 \U14_14_/U2  ( .x(\U14_14_/n2 ), .a(\net222[1] ) );
    inv_1 \U14_14_/U3  ( .x(\U14_14_/n3 ), .a(\net237[1] ) );
    inv_1 \U14_14_/U4  ( .x(\U14_14_/n4 ), .a(\net246[1] ) );
    inv_1 \U14_14_/U5  ( .x(\net212[1] ), .a(\U14_14_/n5 ) );
    and4_1 \U14_15_/U16  ( .x(\U14_15_/n5 ), .a(\U14_15_/n1 ), .b(\U14_15_/n2 
        ), .c(\U14_15_/n3 ), .d(\U14_15_/n4 ) );
    inv_1 \U14_15_/U1  ( .x(\U14_15_/n1 ), .a(\net231[0] ) );
    inv_1 \U14_15_/U2  ( .x(\U14_15_/n2 ), .a(\net222[0] ) );
    inv_1 \U14_15_/U3  ( .x(\U14_15_/n3 ), .a(\net237[0] ) );
    inv_1 \U14_15_/U4  ( .x(\U14_15_/n4 ), .a(\net246[0] ) );
    inv_1 \U14_15_/U5  ( .x(\net212[0] ), .a(\U14_15_/n5 ) );
    and4_1 \U91_0_/U16  ( .x(\U91_0_/n5 ), .a(\U91_0_/n1 ), .b(\U91_0_/n2 ), 
        .c(\U91_0_/n3 ), .d(\U91_0_/n4 ) );
    inv_1 \U91_0_/U1  ( .x(\U91_0_/n1 ), .a(\net219[15] ) );
    inv_1 \U91_0_/U2  ( .x(\U91_0_/n2 ), .a(\net243[15] ) );
    inv_1 \U91_0_/U3  ( .x(\U91_0_/n3 ), .a(\net240[15] ) );
    inv_1 \U91_0_/U4  ( .x(\U91_0_/n4 ), .a(\net228[15] ) );
    inv_1 \U91_0_/U5  ( .x(\net207[15] ), .a(\U91_0_/n5 ) );
    and4_1 \U91_1_/U16  ( .x(\U91_1_/n5 ), .a(\U91_1_/n1 ), .b(\U91_1_/n2 ), 
        .c(\U91_1_/n3 ), .d(\U91_1_/n4 ) );
    inv_1 \U91_1_/U1  ( .x(\U91_1_/n1 ), .a(\net219[14] ) );
    inv_1 \U91_1_/U2  ( .x(\U91_1_/n2 ), .a(\net243[14] ) );
    inv_1 \U91_1_/U3  ( .x(\U91_1_/n3 ), .a(\net240[14] ) );
    inv_1 \U91_1_/U4  ( .x(\U91_1_/n4 ), .a(\net228[14] ) );
    inv_1 \U91_1_/U5  ( .x(\net207[14] ), .a(\U91_1_/n5 ) );
    and4_1 \U91_2_/U16  ( .x(\U91_2_/n5 ), .a(\U91_2_/n1 ), .b(\U91_2_/n2 ), 
        .c(\U91_2_/n3 ), .d(\U91_2_/n4 ) );
    inv_1 \U91_2_/U1  ( .x(\U91_2_/n1 ), .a(\net219[13] ) );
    inv_1 \U91_2_/U2  ( .x(\U91_2_/n2 ), .a(\net243[13] ) );
    inv_1 \U91_2_/U3  ( .x(\U91_2_/n3 ), .a(\net240[13] ) );
    inv_1 \U91_2_/U4  ( .x(\U91_2_/n4 ), .a(\net228[13] ) );
    inv_1 \U91_2_/U5  ( .x(\net207[13] ), .a(\U91_2_/n5 ) );
    and4_1 \U91_3_/U16  ( .x(\U91_3_/n5 ), .a(\U91_3_/n1 ), .b(\U91_3_/n2 ), 
        .c(\U91_3_/n3 ), .d(\U91_3_/n4 ) );
    inv_1 \U91_3_/U1  ( .x(\U91_3_/n1 ), .a(\net219[12] ) );
    inv_1 \U91_3_/U2  ( .x(\U91_3_/n2 ), .a(\net243[12] ) );
    inv_1 \U91_3_/U3  ( .x(\U91_3_/n3 ), .a(\net240[12] ) );
    inv_1 \U91_3_/U4  ( .x(\U91_3_/n4 ), .a(\net228[12] ) );
    inv_1 \U91_3_/U5  ( .x(\net207[12] ), .a(\U91_3_/n5 ) );
    and4_1 \U91_4_/U16  ( .x(\U91_4_/n5 ), .a(\U91_4_/n1 ), .b(\U91_4_/n2 ), 
        .c(\U91_4_/n3 ), .d(\U91_4_/n4 ) );
    inv_1 \U91_4_/U1  ( .x(\U91_4_/n1 ), .a(\net219[11] ) );
    inv_1 \U91_4_/U2  ( .x(\U91_4_/n2 ), .a(\net243[11] ) );
    inv_1 \U91_4_/U3  ( .x(\U91_4_/n3 ), .a(\net240[11] ) );
    inv_1 \U91_4_/U4  ( .x(\U91_4_/n4 ), .a(\net228[11] ) );
    inv_1 \U91_4_/U5  ( .x(\net207[11] ), .a(\U91_4_/n5 ) );
    and4_1 \U91_5_/U16  ( .x(\U91_5_/n5 ), .a(\U91_5_/n1 ), .b(\U91_5_/n2 ), 
        .c(\U91_5_/n3 ), .d(\U91_5_/n4 ) );
    inv_1 \U91_5_/U1  ( .x(\U91_5_/n1 ), .a(\net219[10] ) );
    inv_1 \U91_5_/U2  ( .x(\U91_5_/n2 ), .a(\net243[10] ) );
    inv_1 \U91_5_/U3  ( .x(\U91_5_/n3 ), .a(\net240[10] ) );
    inv_1 \U91_5_/U4  ( .x(\U91_5_/n4 ), .a(\net228[10] ) );
    inv_1 \U91_5_/U5  ( .x(\net207[10] ), .a(\U91_5_/n5 ) );
    and4_1 \U91_6_/U16  ( .x(\U91_6_/n5 ), .a(\U91_6_/n1 ), .b(\U91_6_/n2 ), 
        .c(\U91_6_/n3 ), .d(\U91_6_/n4 ) );
    inv_1 \U91_6_/U1  ( .x(\U91_6_/n1 ), .a(\net219[9] ) );
    inv_1 \U91_6_/U2  ( .x(\U91_6_/n2 ), .a(\net243[9] ) );
    inv_1 \U91_6_/U3  ( .x(\U91_6_/n3 ), .a(\net240[9] ) );
    inv_1 \U91_6_/U4  ( .x(\U91_6_/n4 ), .a(\net228[9] ) );
    inv_1 \U91_6_/U5  ( .x(\net207[9] ), .a(\U91_6_/n5 ) );
    and4_1 \U91_7_/U16  ( .x(\U91_7_/n5 ), .a(\U91_7_/n1 ), .b(\U91_7_/n2 ), 
        .c(\U91_7_/n3 ), .d(\U91_7_/n4 ) );
    inv_1 \U91_7_/U1  ( .x(\U91_7_/n1 ), .a(\net219[8] ) );
    inv_1 \U91_7_/U2  ( .x(\U91_7_/n2 ), .a(\net243[8] ) );
    inv_1 \U91_7_/U3  ( .x(\U91_7_/n3 ), .a(\net240[8] ) );
    inv_1 \U91_7_/U4  ( .x(\U91_7_/n4 ), .a(\net228[8] ) );
    inv_1 \U91_7_/U5  ( .x(\net207[8] ), .a(\U91_7_/n5 ) );
    and4_1 \U91_8_/U16  ( .x(\U91_8_/n5 ), .a(\U91_8_/n1 ), .b(\U91_8_/n2 ), 
        .c(\U91_8_/n3 ), .d(\U91_8_/n4 ) );
    inv_1 \U91_8_/U1  ( .x(\U91_8_/n1 ), .a(\net219[7] ) );
    inv_1 \U91_8_/U2  ( .x(\U91_8_/n2 ), .a(\net243[7] ) );
    inv_1 \U91_8_/U3  ( .x(\U91_8_/n3 ), .a(\net240[7] ) );
    inv_1 \U91_8_/U4  ( .x(\U91_8_/n4 ), .a(\net228[7] ) );
    inv_1 \U91_8_/U5  ( .x(\net207[7] ), .a(\U91_8_/n5 ) );
    and4_1 \U91_9_/U16  ( .x(\U91_9_/n5 ), .a(\U91_9_/n1 ), .b(\U91_9_/n2 ), 
        .c(\U91_9_/n3 ), .d(\U91_9_/n4 ) );
    inv_1 \U91_9_/U1  ( .x(\U91_9_/n1 ), .a(\net219[6] ) );
    inv_1 \U91_9_/U2  ( .x(\U91_9_/n2 ), .a(\net243[6] ) );
    inv_1 \U91_9_/U3  ( .x(\U91_9_/n3 ), .a(\net240[6] ) );
    inv_1 \U91_9_/U4  ( .x(\U91_9_/n4 ), .a(\net228[6] ) );
    inv_1 \U91_9_/U5  ( .x(\net207[6] ), .a(\U91_9_/n5 ) );
    and4_1 \U91_10_/U16  ( .x(\U91_10_/n5 ), .a(\U91_10_/n1 ), .b(\U91_10_/n2 
        ), .c(\U91_10_/n3 ), .d(\U91_10_/n4 ) );
    inv_1 \U91_10_/U1  ( .x(\U91_10_/n1 ), .a(\net219[5] ) );
    inv_1 \U91_10_/U2  ( .x(\U91_10_/n2 ), .a(\net243[5] ) );
    inv_1 \U91_10_/U3  ( .x(\U91_10_/n3 ), .a(\net240[5] ) );
    inv_1 \U91_10_/U4  ( .x(\U91_10_/n4 ), .a(\net228[5] ) );
    inv_1 \U91_10_/U5  ( .x(\net207[5] ), .a(\U91_10_/n5 ) );
    and4_1 \U91_11_/U16  ( .x(\U91_11_/n5 ), .a(\U91_11_/n1 ), .b(\U91_11_/n2 
        ), .c(\U91_11_/n3 ), .d(\U91_11_/n4 ) );
    inv_1 \U91_11_/U1  ( .x(\U91_11_/n1 ), .a(\net219[4] ) );
    inv_1 \U91_11_/U2  ( .x(\U91_11_/n2 ), .a(\net243[4] ) );
    inv_1 \U91_11_/U3  ( .x(\U91_11_/n3 ), .a(\net240[4] ) );
    inv_1 \U91_11_/U4  ( .x(\U91_11_/n4 ), .a(\net228[4] ) );
    inv_1 \U91_11_/U5  ( .x(\net207[4] ), .a(\U91_11_/n5 ) );
    and4_1 \U91_12_/U16  ( .x(\U91_12_/n5 ), .a(\U91_12_/n1 ), .b(\U91_12_/n2 
        ), .c(\U91_12_/n3 ), .d(\U91_12_/n4 ) );
    inv_1 \U91_12_/U1  ( .x(\U91_12_/n1 ), .a(\net219[3] ) );
    inv_1 \U91_12_/U2  ( .x(\U91_12_/n2 ), .a(\net243[3] ) );
    inv_1 \U91_12_/U3  ( .x(\U91_12_/n3 ), .a(\net240[3] ) );
    inv_1 \U91_12_/U4  ( .x(\U91_12_/n4 ), .a(\net228[3] ) );
    inv_1 \U91_12_/U5  ( .x(\net207[3] ), .a(\U91_12_/n5 ) );
    and4_1 \U91_13_/U16  ( .x(\U91_13_/n5 ), .a(\U91_13_/n1 ), .b(\U91_13_/n2 
        ), .c(\U91_13_/n3 ), .d(\U91_13_/n4 ) );
    inv_1 \U91_13_/U1  ( .x(\U91_13_/n1 ), .a(\net219[2] ) );
    inv_1 \U91_13_/U2  ( .x(\U91_13_/n2 ), .a(\net243[2] ) );
    inv_1 \U91_13_/U3  ( .x(\U91_13_/n3 ), .a(\net240[2] ) );
    inv_1 \U91_13_/U4  ( .x(\U91_13_/n4 ), .a(\net228[2] ) );
    inv_1 \U91_13_/U5  ( .x(\net207[2] ), .a(\U91_13_/n5 ) );
    and4_1 \U91_14_/U16  ( .x(\U91_14_/n5 ), .a(\U91_14_/n1 ), .b(\U91_14_/n2 
        ), .c(\U91_14_/n3 ), .d(\U91_14_/n4 ) );
    inv_1 \U91_14_/U1  ( .x(\U91_14_/n1 ), .a(\net219[1] ) );
    inv_1 \U91_14_/U2  ( .x(\U91_14_/n2 ), .a(\net243[1] ) );
    inv_1 \U91_14_/U3  ( .x(\U91_14_/n3 ), .a(\net240[1] ) );
    inv_1 \U91_14_/U4  ( .x(\U91_14_/n4 ), .a(\net228[1] ) );
    inv_1 \U91_14_/U5  ( .x(\net207[1] ), .a(\U91_14_/n5 ) );
    and4_1 \U91_15_/U16  ( .x(\U91_15_/n5 ), .a(\U91_15_/n1 ), .b(\U91_15_/n2 
        ), .c(\U91_15_/n3 ), .d(\U91_15_/n4 ) );
    inv_1 \U91_15_/U1  ( .x(\U91_15_/n1 ), .a(\net219[0] ) );
    inv_1 \U91_15_/U2  ( .x(\U91_15_/n2 ), .a(\net243[0] ) );
    inv_1 \U91_15_/U3  ( .x(\U91_15_/n3 ), .a(\net240[0] ) );
    inv_1 \U91_15_/U4  ( .x(\U91_15_/n4 ), .a(\net228[0] ) );
    inv_1 \U91_15_/U5  ( .x(\net207[0] ), .a(\U91_15_/n5 ) );
    or3_2 \U93_0_/U12  ( .x(chainl[0]), .a(\net207[15] ), .b(\net217[15] ), 
        .c(\net212[15] ) );
    or3_2 \U93_1_/U12  ( .x(chainl[1]), .a(\net207[14] ), .b(\net217[14] ), 
        .c(\net212[14] ) );
    or3_2 \U93_2_/U12  ( .x(chainl[2]), .a(\net207[13] ), .b(\net217[13] ), 
        .c(\net212[13] ) );
    or3_2 \U93_3_/U12  ( .x(chainl[3]), .a(\net207[12] ), .b(\net217[12] ), 
        .c(\net212[12] ) );
    or3_2 \U93_4_/U12  ( .x(chainl[4]), .a(\net207[11] ), .b(\net217[11] ), 
        .c(\net212[11] ) );
    or3_2 \U93_5_/U12  ( .x(chainl[5]), .a(\net207[10] ), .b(\net217[10] ), 
        .c(\net212[10] ) );
    or3_2 \U93_6_/U12  ( .x(chainl[6]), .a(\net207[9] ), .b(\net217[9] ), .c(
        \net212[9] ) );
    or3_2 \U93_7_/U12  ( .x(chainl[7]), .a(\net207[8] ), .b(\net217[8] ), .c(
        \net212[8] ) );
    or3_2 \U93_8_/U12  ( .x(chainh[0]), .a(\net207[7] ), .b(\net217[7] ), .c(
        \net212[7] ) );
    or3_2 \U93_9_/U12  ( .x(chainh[1]), .a(\net207[6] ), .b(\net217[6] ), .c(
        \net212[6] ) );
    or3_2 \U93_10_/U12  ( .x(chainh[2]), .a(\net207[5] ), .b(\net217[5] ), .c(
        \net212[5] ) );
    or3_2 \U93_11_/U12  ( .x(chainh[3]), .a(\net207[4] ), .b(\net217[4] ), .c(
        \net212[4] ) );
    or3_2 \U93_12_/U12  ( .x(chainh[4]), .a(\net207[3] ), .b(\net217[3] ), .c(
        \net212[3] ) );
    or3_2 \U93_13_/U12  ( .x(chainh[5]), .a(\net207[2] ), .b(\net217[2] ), .c(
        \net212[2] ) );
    or3_2 \U93_14_/U12  ( .x(chainh[6]), .a(\net207[1] ), .b(\net217[1] ), .c(
        \net212[1] ) );
    or3_2 \U93_15_/U12  ( .x(chainh[7]), .a(\net207[0] ), .b(\net217[0] ), .c(
        \net212[0] ) );
    inv_1 \U152/U3  ( .x(net198), .a(sendreq) );
    ao23_1 \U158/U19/U21/U1/U1  ( .x(net131), .a(net132), .b(net131), .c(
        net132), .d(rnw[1]), .e(rnw[1]) );
    ao23_1 \U157/U19/U21/U1/U1  ( .x(net176), .a(net132), .b(net176), .c(
        net132), .d(rnw[0]), .e(rnw[0]) );
    ao222_1 \U123/U18/U1/U1  ( .x(net136), .a(net185), .b(net187), .c(net185), 
        .d(net136), .e(net187), .f(net136) );
    aoi21_1 \U151/U30/U1/U1  ( .x(\hdr[4] ), .a(\U151/Z ), .b(net138), .c(
        net198) );
    inv_1 \U151/U30/U1/U2  ( .x(\U151/Z ), .a(\hdr[4] ) );
    nor3_1 \U148/U21/Unr  ( .x(\U148/U21/nr ), .a(net191), .b(net136), .c(
        net293) );
    nand3_1 \U148/U21/Und  ( .x(\U148/U21/nd ), .a(net191), .b(net136), .c(
        net293) );
    oa21_1 \U148/U21/U1  ( .x(\U148/U21/n2 ), .a(\U148/U21/n2 ), .b(
        \U148/U21/nr ), .c(\U148/U21/nd ) );
    inv_1 \U148/U21/U3  ( .x(ack), .a(\U148/U21/n2 ) );
    buf_3 U1 ( .x(n1), .a(net138) );
    buf_3 U2 ( .x(net138), .a(nia) );
    buf_3 U3 ( .x(net269), .a(net146) );
    buf_3 U4 ( .x(net255), .a(\bs[5] ) );
    buf_3 U5 ( .x(net253), .a(\bs[2] ) );
    buf_3 U6 ( .x(net267), .a(\bs[6] ) );
    buf_3 U7 ( .x(net263), .a(\bs[7] ) );
    buf_3 U8 ( .x(net249), .a(\bs[8] ) );
    buf_3 U9 ( .x(net251), .a(\bs[4] ) );
    buf_3 U10 ( .x(net265), .a(\bs[0] ) );
    buf_3 U11 ( .x(net261), .a(\bs[1] ) );
    buf_3 U12 ( .x(net259), .a(\bs[3] ) );
    and2_1 U13 ( .x(\U40_2_/n5 ), .a(\U40_2_/n3 ), .b(\U40_2_/n4 ) );
    and2_1 U14 ( .x(\U40_1_/n5 ), .a(\U40_1_/n3 ), .b(\U40_1_/n4 ) );
    and2_1 U15 ( .x(\U40_9_/n5 ), .a(\U40_9_/n3 ), .b(\U40_9_/n4 ) );
    and2_1 U16 ( .x(\U40_8_/n5 ), .a(\U40_8_/n3 ), .b(\U40_8_/n4 ) );
    and2_1 U17 ( .x(\U40_13_/n5 ), .a(\U40_13_/n3 ), .b(\U40_13_/n4 ) );
    and2_1 U18 ( .x(\U40_0_/n5 ), .a(\U40_0_/n3 ), .b(\U40_0_/n4 ) );
    and2_1 U19 ( .x(\U40_5_/n5 ), .a(\U40_5_/n3 ), .b(\U40_5_/n4 ) );
    and2_1 U20 ( .x(\U40_4_/n5 ), .a(\U40_4_/n3 ), .b(\U40_4_/n4 ) );
    and3_1 U21 ( .x(\U14_12_/n5 ), .a(\U14_12_/n2 ), .b(\U14_12_/n4 ), .c(
        \U14_12_/n1 ) );
    and2_1 U22 ( .x(\U40_12_/n5 ), .a(\U40_12_/n3 ), .b(\U40_12_/n4 ) );
    and2_1 U23 ( .x(\U40_3_/n5 ), .a(\U40_3_/n3 ), .b(\U40_3_/n4 ) );
    and3_1 U24 ( .x(\U14_11_/n5 ), .a(\U14_11_/n2 ), .b(\U14_11_/n4 ), .c(
        \U14_11_/n1 ) );
    and2_1 U25 ( .x(\U40_11_/n5 ), .a(\U40_11_/n3 ), .b(\U40_11_/n4 ) );
    and2_1 U26 ( .x(\U40_10_/n5 ), .a(\U40_10_/n3 ), .b(\U40_10_/n4 ) );
    and2_1 U27 ( .x(\U40_15_/n5 ), .a(\U40_15_/n3 ), .b(\U40_15_/n4 ) );
    and2_1 U28 ( .x(\U40_7_/n5 ), .a(\U40_7_/n3 ), .b(\U40_7_/n4 ) );
    and2_1 U29 ( .x(\U40_6_/n5 ), .a(\U40_6_/n3 ), .b(\U40_6_/n4 ) );
    and2_1 U30 ( .x(\U40_14_/n5 ), .a(\U40_14_/n3 ), .b(\U40_14_/n4 ) );
endmodule


module chain_ic_ctrl_0 ( ack, candefer, eop, nstatack, pltxreq, routetxreq, 
    tok_ack, accept, candefer_ack, defer, eopack, lock, nReset, pltxack, 
    routetxack, tok_err, tok_ok );
input  [1:0] candefer_ack;
input  [1:0] lock;
input  accept, defer, eopack, nReset, pltxack, routetxack, tok_err, tok_ok;
output ack, candefer, eop, nstatack, pltxreq, routetxreq, tok_ack;
    wire \locked[1] , \locked[0] , net21, net12, net20, net16, net10, net7, 
        net6, retry, net27, txnodefer, net13, txunlocked, net5, txmaydefer, 
        txdone, net8, txlocked, net29, net2, net4, lockcleared, net28, net18, 
        net22, net14, net9, net24, net19, net31, net11, net30, net17, net3, 
        reset, net26, nlclear, lwrite, net15, net23, net25, \U249/n5 , 
        \U249/n1 , \U249/n2 , \U249/n3 , \U249/n4 , \U286/U28/U1/clr , 
        \U286/U28/U1/set , \U285/U28/U1/clr , \U285/U28/U1/set , 
        \U262/U25/U1/clr , \U262/U25/U1/ob , \U284/U25/U1/clr , 
        \U284/U25/U1/ob , \U283/U25/U1/clr , \U283/U25/U1/ob , \U288/Z , 
        \U289/Z , \U287/Z , \U149/nr , \U149/nd , \U149/n2 , \U160/acb , 
        \U160/U1/Z , \U136/nlsense , \U136/nulsense , \U136/nwh , \U136/nwl , 
        \U136/nclear_latch , n1, n2;
    nand2_1 \U146/U5  ( .x(candefer), .a(net23), .b(net25) );
    or2_1 \U277/U12  ( .x(net6), .a(net19), .b(net9) );
    or2_1 \U264/U12  ( .x(retry), .a(net31), .b(net24) );
    or2_1 \U259/U12  ( .x(net28), .a(net27), .b(net7) );
    or2_1 \U140/U12  ( .x(net18), .a(net13), .b(net8) );
    or2_1 \U148/U12  ( .x(net11), .a(net15), .b(routetxack) );
    and4_1 \U249/U16  ( .x(\U249/n5 ), .a(\U249/n1 ), .b(\U249/n2 ), .c(
        \U249/n3 ), .d(\U249/n4 ) );
    inv_1 \U249/U1  ( .x(\U249/n1 ), .a(txnodefer) );
    inv_1 \U249/U2  ( .x(\U249/n2 ), .a(net16) );
    inv_1 \U249/U3  ( .x(\U249/n3 ), .a(net9) );
    inv_1 \U249/U4  ( .x(\U249/n4 ), .a(net19) );
    inv_1 \U249/U5  ( .x(ack), .a(\U249/n5 ) );
    nor3_2 \U40/U16  ( .x(nstatack), .a(net16), .b(reset), .c(retry) );
    nor3_2 \U275/U16  ( .x(net17), .a(net29), .b(reset), .c(tok_ack) );
    buf_3 \U290/U8  ( .x(net12), .a(txmaydefer) );
    nor2_1 \U154/U5  ( .x(nlclear), .a(net4), .b(net31) );
    or2_2 \U274/U12  ( .x(pltxreq), .a(net22), .b(net14) );
    or3_1 \U260/U12  ( .x(eop), .a(net31), .b(txlocked), .c(net4) );
    inv_1 \U147/U3  ( .x(net3), .a(net29) );
    inv_1 \U174/U3  ( .x(reset), .a(nReset) );
    aoai211_1 \U286/U28/U1/U1  ( .x(\U286/U28/U1/clr ), .a(net3), .b(n1), .c(
        net17), .d(net22) );
    nand3_1 \U286/U28/U1/U2  ( .x(\U286/U28/U1/set ), .a(net17), .b(net3), .c(
        n1) );
    nand2_2 \U286/U28/U1/U3  ( .x(net22), .a(\U286/U28/U1/clr ), .b(
        \U286/U28/U1/set ) );
    aoai211_1 \U285/U28/U1/U1  ( .x(\U285/U28/U1/clr ), .a(net3), .b(n2), .c(
        net17), .d(net14) );
    nand3_1 \U285/U28/U1/U2  ( .x(\U285/U28/U1/set ), .a(net17), .b(net3), .c(
        n2) );
    nand2_2 \U285/U28/U1/U3  ( .x(net14), .a(\U285/U28/U1/clr ), .b(
        \U285/U28/U1/set ) );
    ao222_1 \U254/U18/U1/U1  ( .x(net31), .a(defer), .b(txunlocked), .c(defer), 
        .d(net31), .e(txunlocked), .f(net31) );
    ao222_1 \U252/U18/U1/U1  ( .x(net19), .a(tok_err), .b(net12), .c(tok_err), 
        .d(net19), .e(net12), .f(net19) );
    ao222_1 \U276/U18/U1/U1  ( .x(net24), .a(txlocked), .b(defer), .c(txlocked
        ), .d(net24), .e(defer), .f(net24) );
    ao222_1 \U251/U18/U1/U1  ( .x(net9), .a(tok_ok), .b(net12), .c(tok_ok), 
        .d(net9), .e(net12), .f(net9) );
    ao222_1 \U235/U18/U1/U1  ( .x(tok_ack), .a(ack), .b(net2), .c(ack), .d(
        tok_ack), .e(net2), .f(tok_ack) );
    ao222_1 \U247/U18/U1/U1  ( .x(txnodefer), .a(txdone), .b(candefer_ack[0]), 
        .c(txdone), .d(txnodefer), .e(candefer_ack[0]), .f(txnodefer) );
    ao222_2 \U246/U19/U1/U1  ( .x(txlocked), .a(net14), .b(txdone), .c(net14), 
        .d(txlocked), .e(txdone), .f(txlocked) );
    ao222_2 \U245/U19/U1/U1  ( .x(txunlocked), .a(txdone), .b(net22), .c(
        txdone), .d(txunlocked), .e(net22), .f(txunlocked) );
    ao222_1 \U269/U18/U1/U1  ( .x(net2), .a(net28), .b(net18), .c(net28), .d(
        net2), .e(net18), .f(net2) );
    ao222_1 \U268/U18/U1/U1  ( .x(net5), .a(eopack), .b(lockcleared), .c(
        eopack), .d(net5), .e(lockcleared), .f(net5) );
    ao222_1 \U256/U18/U1/U1  ( .x(net4), .a(tok_err), .b(txunlocked), .c(
        tok_err), .d(net4), .e(txunlocked), .f(net4) );
    ao222_1 \U175/U18/U1/U1  ( .x(net29), .a(net2), .b(retry), .c(net2), .d(
        net29), .e(retry), .f(net29) );
    ao222_1 \U255/U18/U1/U1  ( .x(net8), .a(txlocked), .b(eopack), .c(txlocked
        ), .d(net8), .e(eopack), .f(net8) );
    ao222_2 \U248/U19/U1/U1  ( .x(txmaydefer), .a(candefer_ack[1]), .b(txdone), 
        .c(candefer_ack[1]), .d(txmaydefer), .e(txdone), .f(txmaydefer) );
    ao222_2 \U250/U19/U1/U1  ( .x(net16), .a(accept), .b(net12), .c(accept), 
        .d(net16), .e(net12), .f(net16) );
    oa31_1 \U262/U25/U1/Uclr  ( .x(\U262/U25/U1/clr ), .a(txunlocked), .b(net5
        ), .c(tok_ok), .d(net13) );
    oaoi211_1 \U262/U25/U1/Uaoi  ( .x(\U262/U25/U1/ob ), .a(net5), .b(tok_ok), 
        .c(txunlocked), .d(\U262/U25/U1/clr ) );
    inv_2 \U262/U25/U1/Ui  ( .x(net13), .a(\U262/U25/U1/ob ) );
    oa31_1 \U284/U25/U1/Uclr  ( .x(\U284/U25/U1/clr ), .a(txnodefer), .b(
        tok_ok), .c(tok_err), .d(net27) );
    oaoi211_1 \U284/U25/U1/Uaoi  ( .x(\U284/U25/U1/ob ), .a(tok_ok), .b(
        tok_err), .c(txnodefer), .d(\U284/U25/U1/clr ) );
    inv_2 \U284/U25/U1/Ui  ( .x(net27), .a(\U284/U25/U1/ob ) );
    oa31_1 \U283/U25/U1/Uclr  ( .x(\U283/U25/U1/clr ), .a(net10), .b(net6), 
        .c(retry), .d(net7) );
    oaoi211_1 \U283/U25/U1/Uaoi  ( .x(\U283/U25/U1/ob ), .a(net6), .b(retry), 
        .c(net10), .d(\U283/U25/U1/clr ) );
    inv_2 \U283/U25/U1/Ui  ( .x(net7), .a(\U283/U25/U1/ob ) );
    aoi21_1 \U289/U30/U1/U1  ( .x(net20), .a(\U289/Z ), .b(net16), .c(net12)
         );
    inv_1 \U289/U30/U1/U2  ( .x(\U289/Z ), .a(net20) );
    aoi21_1 \U287/U30/U1/U1  ( .x(net21), .a(\U287/Z ), .b(accept), .c(net12)
         );
    inv_1 \U287/U30/U1/U2  ( .x(\U287/Z ), .a(net21) );
    aoi222_1 \U288/U30/U1  ( .x(net10), .a(net20), .b(net21), .c(net20), .d(
        \U288/Z ), .e(net21), .f(\U288/Z ) );
    inv_1 \U288/U30/Uinv  ( .x(\U288/Z ), .a(net10) );
    nor3_1 \U149/Unr  ( .x(\U149/nr ), .a(pltxack), .b(net11), .c(net30) );
    nand3_1 \U149/Und  ( .x(\U149/nd ), .a(pltxack), .b(net11), .c(net30) );
    oa21_1 \U149/U1  ( .x(\U149/n2 ), .a(\U149/n2 ), .b(\U149/nr ), .c(
        \U149/nd ) );
    inv_2 \U149/U3  ( .x(txdone), .a(\U149/n2 ) );
    inv_1 \U133/U618/U3  ( .x(net23), .a(net15) );
    inv_1 \U133/U617/U3  ( .x(net25), .a(routetxreq) );
    ao23_1 \U133/U616/U21/U1/U1  ( .x(routetxreq), .a(pltxreq), .b(routetxreq), 
        .c(pltxreq), .d(\locked[0] ), .e(net23) );
    ao23_1 \U133/U615/U21/U1/U1  ( .x(net15), .a(pltxreq), .b(net15), .c(
        pltxreq), .d(\locked[1] ), .e(net25) );
    and2_1 \U160/U2/U8  ( .x(lwrite), .a(candefer), .b(\U160/acb ) );
    nor2_1 \U160/U3/U5  ( .x(net30), .a(\U160/acb ), .b(net26) );
    oai21_1 \U160/U1/U30/U1/U1  ( .x(\U160/acb ), .a(\U160/U1/Z ), .b(net26), 
        .c(candefer) );
    inv_1 \U160/U1/U30/U1/U2  ( .x(\U160/U1/Z ), .a(\U160/acb ) );
    nand3_2 \U136/U48/U16  ( .x(\locked[0] ), .a(\locked[1] ), .b(
        \U136/nclear_latch ), .c(\U136/nwl ) );
    nor2_0 \U136/U36/U5  ( .x(\U136/nulsense ), .a(\locked[1] ), .b(\U136/nwl 
        ) );
    nor2_0 \U136/U37/U5  ( .x(\U136/nlsense ), .a(\U136/nwh ), .b(\locked[0] )
         );
    and2_1 \U136/U76/U8  ( .x(\U136/nclear_latch ), .a(nReset), .b(nlclear) );
    nor2_1 \U136/U77/U5  ( .x(lockcleared), .a(nlclear), .b(\locked[1] ) );
    nand2_1 \U136/U14/U5  ( .x(\U136/nwl ), .a(lwrite), .b(n2) );
    nand2_1 \U136/U15/U5  ( .x(\U136/nwh ), .a(n1), .b(lwrite) );
    nand2_2 \U136/U47/U5  ( .x(\locked[1] ), .a(\U136/nwh ), .b(\locked[0] )
         );
    or2_4 \U136/U35/U12  ( .x(net26), .a(\U136/nlsense ), .b(\U136/nulsense )
         );
    buf_1 U1 ( .x(n1), .a(lock[1]) );
    buf_1 U2 ( .x(n2), .a(lock[0]) );
endmodule


module chain_irdemuxNew_0 ( err, ncback, rd, rnw, status, cbh, cbl, nReset, 
    nack, statusack );
output [1:0] err;
output [63:0] rd;
output [1:0] rnw;
output [1:0] status;
input  [7:0] cbh;
input  [7:0] cbl;
input  nReset, nack, statusack;
output ncback;
    wire n17, n18, \ncd[7] , \ncd[6] , \ncd[5] , \ncd[4] , \ncd[3] , \ncd[2] , 
        \ncd[1] , \ncd[0] , \col_h[2] , \col_h[1] , \col_h[0] , \col_l[2] , 
        \col_l[1] , \col_l[0] , \opc_l[2] , \opc_l[1] , \opc_l[0] , \opc_h[1] , 
        \opc_h[0] , pullcd, net86, net171, net168, net103, net170, bpullcd, 
        reset, net94, read_lhw, net166, net169, read, net139, net172, 
        start_receiving, net193, net167, net149, net173, pkt_normal, notify, 
        net150, write, net176, net162, pkt_done, net0187, net0208, 
        \U1697/U21/nr , \U1697/U21/nd , \U1697/U21/n2 , \U307/U21/nr , 
        \U307/U21/nd , \U307/U21/n2 , \U1664/U28/Z , \U1664/U32/Z , 
        \U1664/U29/Z , \U1664/U33/Z , \U1664/U30/Z , \U1664/U31/Z , 
        \U1664/U37/Z , \U1664/y[0] , \U1664/y[1] , \U1664/x[1] , \U1664/x[3] , 
        \U1664/x[2] , \U1664/x[0] , \U1698/nr , \U1698/nd , \U1698/n2 , 
        \I6/oh[7] , \I6/oh[6] , \I6/oh[4] , \I6/oh[3] , \I6/oh[2] , \I6/ol[7] , 
        \I6/ol[6] , \I6/ol[4] , \I6/ol[3] , \I6/drivel , \I6/driveh , 
        \I6/localcd , \I6/ncd[7] , \I6/ncd[6] , \I6/ncd[5] , \I6/ncd[4] , 
        \I6/ncd[3] , \I6/ncd[2] , \I6/ncd[1] , \I6/ncd[0] , \I6/ba , 
        \I6/latch , \I6/acb , \I6/ctrlack_internal , \I6/nlocalcd , 
        \I6/U4/U28/U1/clr , \I6/U4/U28/U1/set , \I6/U1/Z , \I6/U1664/y[0] , 
        \I6/U1664/y[1] , \I6/U1664/x[1] , \I6/U1664/x[3] , \I6/U1664/x[2] , 
        \I6/U1664/x[0] , \I6/U1664/U28/Z , \I6/U1664/U32/Z , \I6/U1664/U29/Z , 
        \I6/U1664/U33/Z , \I6/U1664/U30/Z , \I6/U1664/U31/Z , \I6/U1664/U37/Z , 
        \I6/U1669/nr , \I6/U1669/nd , \I6/U1669/n2 , \U1667/drivel , 
        \U1667/driveh , \U1667/localcd , \U1667/ncd[7] , \U1667/ncd[6] , 
        \U1667/ncd[5] , \U1667/ncd[4] , \U1667/ncd[3] , \U1667/ncd[2] , 
        \U1667/ncd[1] , \U1667/ncd[0] , \U1667/ba , \U1667/latch , \U1667/acb , 
        \U1667/ctrlack_internal , \U1667/nlocalcd , \U1667/U4/U28/U1/clr , 
        \U1667/U4/U28/U1/set , \U1667/U1/Z , \U1667/U1664/y[0] , 
        \U1667/U1664/y[1] , \U1667/U1664/x[1] , \U1667/U1664/x[3] , 
        \U1667/U1664/x[2] , \U1667/U1664/x[0] , \U1667/U1664/U28/Z , 
        \U1667/U1664/U32/Z , \U1667/U1664/U29/Z , \U1667/U1664/U33/Z , 
        \U1667/U1664/U30/Z , \U1667/U1664/U31/Z , \U1667/U1664/U37/Z , 
        \U1667/U1669/nr , \U1667/U1669/nd , \U1667/U1669/n2 , \U1650/oh[4] , 
        \U1650/oh[3] , \U1650/oh[2] , \U1650/oh[1] , \U1650/oh[0] , 
        \U1650/ol[4] , \U1650/ol[3] , \U1650/ol[2] , \U1650/ol[1] , 
        \U1650/ol[0] , \U1650/drivel , \U1650/driveh , \U1650/localcd , 
        \U1650/ncd[7] , \U1650/ncd[6] , \U1650/ncd[5] , \U1650/ncd[4] , 
        \U1650/ncd[3] , \U1650/ncd[2] , \U1650/ncd[1] , \U1650/ncd[0] , 
        \U1650/ba , \U1650/latch , \U1650/acb , \U1650/ctrlack_internal , 
        \U1650/nlocalcd , \U1650/U4/U28/U1/clr , \U1650/U4/U28/U1/set , 
        \U1650/U1/Z , \U1650/U1664/y[0] , \U1650/U1664/y[1] , 
        \U1650/U1664/x[1] , \U1650/U1664/x[3] , \U1650/U1664/x[2] , 
        \U1650/U1664/x[0] , \U1650/U1664/U28/Z , \U1650/U1664/U32/Z , 
        \U1650/U1664/U29/Z , \U1650/U1664/U33/Z , \U1650/U1664/U30/Z , 
        \U1650/U1664/U31/Z , \U1650/U1664/U37/Z , \U1650/U1669/nr , 
        \U1650/U1669/nd , \U1650/U1669/n2 , \U1666/drivel , \U1666/driveh , 
        \U1666/localcd , \U1666/ncd[7] , \U1666/ncd[6] , \U1666/ncd[5] , 
        \U1666/ncd[4] , \U1666/ncd[3] , \U1666/ncd[2] , \U1666/ncd[1] , 
        \U1666/ncd[0] , \U1666/ba , \U1666/latch , \U1666/acb , 
        \U1666/ctrlack_internal , \U1666/nlocalcd , \U1666/U4/U28/U1/clr , 
        \U1666/U4/U28/U1/set , \U1666/U1/Z , \U1666/U1664/y[0] , 
        \U1666/U1664/y[1] , \U1666/U1664/x[1] , \U1666/U1664/x[3] , 
        \U1666/U1664/x[2] , \U1666/U1664/x[0] , \U1666/U1664/U28/Z , 
        \U1666/U1664/U32/Z , \U1666/U1664/U29/Z , \U1666/U1664/U33/Z , 
        \U1666/U1664/U30/Z , \U1666/U1664/U31/Z , \U1666/U1664/U37/Z , 
        \U1666/U1669/nr , \U1666/U1669/nd , \U1666/U1669/n2 , \I1/drivel , 
        \I1/driveh , \I1/localcd , \I1/ncd[7] , \I1/ncd[6] , \I1/ncd[5] , 
        \I1/ncd[4] , \I1/ncd[3] , \I1/ncd[2] , \I1/ncd[1] , \I1/ncd[0] , 
        \I1/ba , \I1/latch , \I1/acb , \I1/ctrlack_internal , \I1/nlocalcd , 
        \I1/U4/U28/U1/clr , \I1/U4/U28/U1/set , \I1/U1/Z , \I1/U1664/y[0] , 
        \I1/U1664/y[1] , \I1/U1664/x[1] , \I1/U1664/x[3] , \I1/U1664/x[2] , 
        \I1/U1664/x[0] , \I1/U1664/U28/Z , \I1/U1664/U32/Z , \I1/U1664/U29/Z , 
        \I1/U1664/U33/Z , \I1/U1664/U30/Z , \I1/U1664/U31/Z , \I1/U1664/U37/Z , 
        \I1/U1669/nr , \I1/U1669/nd , \I1/U1669/n2 , \I2/drivel , \I2/driveh , 
        \I2/localcd , \I2/ncd[7] , \I2/ncd[6] , \I2/ncd[5] , \I2/ncd[4] , 
        \I2/ncd[3] , \I2/ncd[2] , \I2/ncd[1] , \I2/ncd[0] , \I2/ba , 
        \I2/latch , \I2/acb , \I2/ctrlack_internal , \I2/nlocalcd , 
        \I2/U4/U28/U1/clr , \I2/U4/U28/U1/set , \I2/U1/Z , \I2/U1664/y[0] , 
        \I2/U1664/y[1] , \I2/U1664/x[1] , \I2/U1664/x[3] , \I2/U1664/x[2] , 
        \I2/U1664/x[0] , \I2/U1664/U28/Z , \I2/U1664/U32/Z , \I2/U1664/U29/Z , 
        \I2/U1664/U33/Z , \I2/U1664/U30/Z , \I2/U1664/U31/Z , \I2/U1664/U37/Z , 
        \I2/U1669/nr , \I2/U1669/nd , \I2/U1669/n2 , n1, n2, n3, n4, n5, n6, 
        n7, n8, n9, n10, n11, n12, n13, n14;
    buf_1 U262 ( .x(bpullcd), .a(pullcd) );
    or2_4 \U1674/U12  ( .x(net162), .a(nack), .b(reset) );
    and2_4 \U1785/U8  ( .x(pkt_normal), .a(\opc_l[2] ), .b(\opc_l[1] ) );
    and2_4 \U1777/U8  ( .x(net150), .a(\opc_l[2] ), .b(\opc_h[1] ) );
    or3_1 \U1813/U12  ( .x(pkt_done), .a(write), .b(reset), .c(net193) );
    nor2_1 \U1651_0_/U5  ( .x(\ncd[0] ), .a(cbh[0]), .b(cbl[0]) );
    nor2_1 \U1651_1_/U5  ( .x(\ncd[1] ), .a(cbh[1]), .b(cbl[1]) );
    nor2_1 \U1651_2_/U5  ( .x(\ncd[2] ), .a(cbh[2]), .b(cbl[2]) );
    nor2_1 \U1651_3_/U5  ( .x(\ncd[3] ), .a(cbh[3]), .b(cbl[3]) );
    nor2_1 \U1651_4_/U5  ( .x(\ncd[4] ), .a(cbh[4]), .b(cbl[4]) );
    nor2_1 \U1651_5_/U5  ( .x(\ncd[5] ), .a(cbh[5]), .b(cbl[5]) );
    nor2_1 \U1651_6_/U5  ( .x(\ncd[6] ), .a(cbh[6]), .b(cbl[6]) );
    nor2_1 \U1651_7_/U5  ( .x(\ncd[7] ), .a(cbh[7]), .b(cbl[7]) );
    nor2_1 \U1812/U5  ( .x(start_receiving), .a(notify), .b(net176) );
    nor2_1 \I7/U5  ( .x(net86), .a(net172), .b(net173) );
    nor2_1 \I4/U5  ( .x(net171), .a(net169), .b(net170) );
    nor2_1 \I3/U5  ( .x(net168), .a(net166), .b(net167) );
    inv_2 \U1675/U3  ( .x(reset), .a(nReset) );
    nand3_2 \U193/U16  ( .x(ncback), .a(net86), .b(net171), .c(net168) );
    ao222_1 \U1811/U18/U1/U1  ( .x(net176), .a(net162), .b(pkt_done), .c(
        net162), .d(net176), .e(pkt_done), .f(net176) );
    aoi222_1 \U1664/U28/U30/U1  ( .x(\U1664/x[3] ), .a(\ncd[7] ), .b(\ncd[6] ), 
        .c(\ncd[7] ), .d(\U1664/U28/Z ), .e(\ncd[6] ), .f(\U1664/U28/Z ) );
    inv_1 \U1664/U28/U30/Uinv  ( .x(\U1664/U28/Z ), .a(\U1664/x[3] ) );
    aoi222_1 \U1664/U32/U30/U1  ( .x(\U1664/x[0] ), .a(\ncd[1] ), .b(\ncd[0] ), 
        .c(\ncd[1] ), .d(\U1664/U32/Z ), .e(\ncd[0] ), .f(\U1664/U32/Z ) );
    inv_1 \U1664/U32/U30/Uinv  ( .x(\U1664/U32/Z ), .a(\U1664/x[0] ) );
    aoi222_1 \U1664/U29/U30/U1  ( .x(\U1664/x[2] ), .a(\ncd[5] ), .b(\ncd[4] ), 
        .c(\ncd[5] ), .d(\U1664/U29/Z ), .e(\ncd[4] ), .f(\U1664/U29/Z ) );
    inv_1 \U1664/U29/U30/Uinv  ( .x(\U1664/U29/Z ), .a(\U1664/x[2] ) );
    aoi222_1 \U1664/U33/U30/U1  ( .x(\U1664/y[0] ), .a(\U1664/x[1] ), .b(
        \U1664/x[0] ), .c(\U1664/x[1] ), .d(\U1664/U33/Z ), .e(\U1664/x[0] ), 
        .f(\U1664/U33/Z ) );
    inv_1 \U1664/U33/U30/Uinv  ( .x(\U1664/U33/Z ), .a(\U1664/y[0] ) );
    aoi222_1 \U1664/U30/U30/U1  ( .x(\U1664/y[1] ), .a(\U1664/x[3] ), .b(
        \U1664/x[2] ), .c(\U1664/x[3] ), .d(\U1664/U30/Z ), .e(\U1664/x[2] ), 
        .f(\U1664/U30/Z ) );
    inv_1 \U1664/U30/U30/Uinv  ( .x(\U1664/U30/Z ), .a(\U1664/y[1] ) );
    aoi222_1 \U1664/U31/U30/U1  ( .x(\U1664/x[1] ), .a(\ncd[3] ), .b(\ncd[2] ), 
        .c(\ncd[3] ), .d(\U1664/U31/Z ), .e(\ncd[2] ), .f(\U1664/U31/Z ) );
    inv_1 \U1664/U31/U30/Uinv  ( .x(\U1664/U31/Z ), .a(\U1664/x[1] ) );
    aoi222_1 \U1664/U37/U30/U1  ( .x(pullcd), .a(\U1664/y[0] ), .b(
        \U1664/y[1] ), .c(\U1664/y[0] ), .d(\U1664/U37/Z ), .e(\U1664/y[1] ), 
        .f(\U1664/U37/Z ) );
    inv_1 \U1664/U37/U30/Uinv  ( .x(\U1664/U37/Z ), .a(pullcd) );
    nor3_1 \U1697/U21/Unr  ( .x(\U1697/U21/nr ), .a(rnw[0]), .b(pkt_normal), 
        .c(net149) );
    nand3_1 \U1697/U21/Und  ( .x(\U1697/U21/nd ), .a(rnw[0]), .b(pkt_normal), 
        .c(net149) );
    oa21_1 \U1697/U21/U1  ( .x(\U1697/U21/n2 ), .a(\U1697/U21/n2 ), .b(
        \U1697/U21/nr ), .c(\U1697/U21/nd ) );
    inv_1 \U1697/U21/U3  ( .x(write), .a(\U1697/U21/n2 ) );
    nor3_1 \U307/U21/Unr  ( .x(\U307/U21/nr ), .a(net149), .b(net150), .c(
        statusack) );
    nand3_1 \U307/U21/Und  ( .x(\U307/U21/nd ), .a(net149), .b(net150), .c(
        statusack) );
    oa21_1 \U307/U21/U1  ( .x(\U307/U21/n2 ), .a(\U307/U21/n2 ), .b(
        \U307/U21/nr ), .c(\U307/U21/nd ) );
    inv_1 \U307/U21/U3  ( .x(notify), .a(\U307/U21/n2 ) );
    nor3_1 \U1698/Unr  ( .x(\U1698/nr ), .a(rnw[1]), .b(pkt_normal), .c(net149
        ) );
    nand3_1 \U1698/Und  ( .x(\U1698/nd ), .a(rnw[1]), .b(pkt_normal), .c(
        net149) );
    oa21_1 \U1698/U1  ( .x(\U1698/n2 ), .a(\U1698/n2 ), .b(\U1698/nr ), .c(
        \U1698/nd ) );
    inv_2 \U1698/U3  ( .x(read), .a(\U1698/n2 ) );
    and2_1 \U1756/U1754/U8  ( .x(n17), .a(\opc_h[0] ), .b(pkt_normal) );
    and2_1 \U1756/U1755/U8  ( .x(n18), .a(\opc_l[0] ), .b(pkt_normal) );
    and2_1 \U1800/U1754/U8  ( .x(rnw[1]), .a(net0187), .b(pkt_normal) );
    and2_1 \U1800/U1755/U8  ( .x(rnw[0]), .a(net0208), .b(pkt_normal) );
    and2_1 \U1758/U1754/U8  ( .x(status[1]), .a(\opc_h[0] ), .b(net150) );
    and2_1 \U1758/U1755/U8  ( .x(status[0]), .a(\opc_l[0] ), .b(net150) );
    buf_2 \I6/U1653  ( .x(\I6/latch ), .a(net173) );
    nor2_1 \I6/U264/U5  ( .x(\I6/nlocalcd ), .a(reset), .b(\I6/localcd ) );
    nor2_1 \I6/U1659_0_/U5  ( .x(\I6/ncd[0] ), .a(\opc_l[0] ), .b(\opc_h[0] )
         );
    nor2_1 \I6/U1659_1_/U5  ( .x(\I6/ncd[1] ), .a(\opc_l[1] ), .b(\opc_h[1] )
         );
    nor2_1 \I6/U1659_2_/U5  ( .x(\I6/ncd[2] ), .a(\opc_l[2] ), .b(\I6/oh[2] )
         );
    nor2_1 \I6/U1659_3_/U5  ( .x(\I6/ncd[3] ), .a(\I6/ol[3] ), .b(\I6/oh[3] )
         );
    nor2_1 \I6/U1659_4_/U5  ( .x(\I6/ncd[4] ), .a(\I6/ol[4] ), .b(\I6/oh[4] )
         );
    nor2_1 \I6/U1659_5_/U5  ( .x(\I6/ncd[5] ), .a(net0208), .b(net0187) );
    nor2_1 \I6/U1659_6_/U5  ( .x(\I6/ncd[6] ), .a(\I6/ol[6] ), .b(\I6/oh[6] )
         );
    nor2_1 \I6/U1659_7_/U5  ( .x(\I6/ncd[7] ), .a(\I6/ol[7] ), .b(\I6/oh[7] )
         );
    nor2_1 \I6/U3/U5  ( .x(\I6/ctrlack_internal ), .a(\I6/acb ), .b(\I6/ba )
         );
    buf_2 \I6/U1665/U7  ( .x(\I6/driveh ), .a(net139) );
    buf_2 \I6/U1666/U7  ( .x(\I6/drivel ), .a(net139) );
    ao23_1 \I6/U1658_0_/U21/U1/U1  ( .x(\opc_l[0] ), .a(\I6/driveh ), .b(
        \opc_l[0] ), .c(\I6/driveh ), .d(cbl[0]), .e(n12) );
    ao23_1 \I6/U1658_1_/U21/U1/U1  ( .x(\opc_l[1] ), .a(\I6/driveh ), .b(
        \opc_l[1] ), .c(\I6/drivel ), .d(cbl[1]), .e(n12) );
    ao23_1 \I6/U1658_2_/U21/U1/U1  ( .x(\opc_l[2] ), .a(\I6/drivel ), .b(
        \opc_l[2] ), .c(n13), .d(cbl[2]), .e(n12) );
    ao23_1 \I6/U1658_3_/U21/U1/U1  ( .x(\I6/ol[3] ), .a(\I6/drivel ), .b(
        \I6/ol[3] ), .c(\I6/drivel ), .d(cbl[3]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_4_/U21/U1/U1  ( .x(\I6/ol[4] ), .a(n13), .b(\I6/ol[4] ), 
        .c(n13), .d(cbl[4]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_5_/U21/U1/U1  ( .x(net0208), .a(\I6/driveh ), .b(net0208), 
        .c(\I6/driveh ), .d(cbl[5]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_6_/U21/U1/U1  ( .x(\I6/ol[6] ), .a(n13), .b(\I6/ol[6] ), 
        .c(n13), .d(cbl[6]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_7_/U21/U1/U1  ( .x(\I6/ol[7] ), .a(n13), .b(\I6/ol[7] ), 
        .c(\I6/driveh ), .d(cbl[7]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_0_/U21/U1/U1  ( .x(\opc_h[0] ), .a(n13), .b(\opc_h[0] ), 
        .c(\I6/drivel ), .d(cbh[0]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_1_/U21/U1/U1  ( .x(\opc_h[1] ), .a(\I6/driveh ), .b(
        \opc_h[1] ), .c(n13), .d(cbh[1]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_2_/U21/U1/U1  ( .x(\I6/oh[2] ), .a(\I6/driveh ), .b(
        \I6/oh[2] ), .c(n13), .d(cbh[2]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_3_/U21/U1/U1  ( .x(\I6/oh[3] ), .a(\I6/drivel ), .b(
        \I6/oh[3] ), .c(\I6/drivel ), .d(cbh[3]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_4_/U21/U1/U1  ( .x(\I6/oh[4] ), .a(n13), .b(\I6/oh[4] ), 
        .c(\I6/driveh ), .d(cbh[4]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_5_/U21/U1/U1  ( .x(net0187), .a(\I6/driveh ), .b(net0187), 
        .c(\I6/driveh ), .d(cbh[5]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_6_/U21/U1/U1  ( .x(\I6/oh[6] ), .a(\I6/drivel ), .b(
        \I6/oh[6] ), .c(\I6/drivel ), .d(cbh[6]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_7_/U21/U1/U1  ( .x(\I6/oh[7] ), .a(\I6/drivel ), .b(
        \I6/oh[7] ), .c(n13), .d(cbh[7]), .e(\I6/latch ) );
    aoai211_1 \I6/U4/U28/U1/U1  ( .x(\I6/U4/U28/U1/clr ), .a(net139), .b(
        \I6/acb ), .c(\I6/nlocalcd ), .d(net173) );
    nand3_1 \I6/U4/U28/U1/U2  ( .x(\I6/U4/U28/U1/set ), .a(\I6/nlocalcd ), .b(
        net139), .c(\I6/acb ) );
    nand2_2 \I6/U4/U28/U1/U3  ( .x(net173), .a(\I6/U4/U28/U1/clr ), .b(
        \I6/U4/U28/U1/set ) );
    oai21_1 \I6/U1/U30/U1/U1  ( .x(\I6/acb ), .a(\I6/U1/Z ), .b(\I6/ba ), .c(
        net139) );
    inv_1 \I6/U1/U30/U1/U2  ( .x(\I6/U1/Z ), .a(\I6/acb ) );
    ao222_1 \I6/U5/U18/U1/U1  ( .x(\I6/ba ), .a(\I6/latch ), .b(n14), .c(
        \I6/latch ), .d(\I6/ba ), .e(n14), .f(\I6/ba ) );
    aoi222_1 \I6/U1664/U28/U30/U1  ( .x(\I6/U1664/x[3] ), .a(\I6/ncd[7] ), .b(
        \I6/ncd[6] ), .c(\I6/ncd[7] ), .d(\I6/U1664/U28/Z ), .e(\I6/ncd[6] ), 
        .f(\I6/U1664/U28/Z ) );
    inv_1 \I6/U1664/U28/U30/Uinv  ( .x(\I6/U1664/U28/Z ), .a(\I6/U1664/x[3] )
         );
    aoi222_1 \I6/U1664/U32/U30/U1  ( .x(\I6/U1664/x[0] ), .a(\I6/ncd[1] ), .b(
        \I6/ncd[0] ), .c(\I6/ncd[1] ), .d(\I6/U1664/U32/Z ), .e(\I6/ncd[0] ), 
        .f(\I6/U1664/U32/Z ) );
    inv_1 \I6/U1664/U32/U30/Uinv  ( .x(\I6/U1664/U32/Z ), .a(\I6/U1664/x[0] )
         );
    aoi222_1 \I6/U1664/U29/U30/U1  ( .x(\I6/U1664/x[2] ), .a(\I6/ncd[5] ), .b(
        \I6/ncd[4] ), .c(\I6/ncd[5] ), .d(\I6/U1664/U29/Z ), .e(\I6/ncd[4] ), 
        .f(\I6/U1664/U29/Z ) );
    inv_1 \I6/U1664/U29/U30/Uinv  ( .x(\I6/U1664/U29/Z ), .a(\I6/U1664/x[2] )
         );
    aoi222_1 \I6/U1664/U33/U30/U1  ( .x(\I6/U1664/y[0] ), .a(\I6/U1664/x[1] ), 
        .b(\I6/U1664/x[0] ), .c(\I6/U1664/x[1] ), .d(\I6/U1664/U33/Z ), .e(
        \I6/U1664/x[0] ), .f(\I6/U1664/U33/Z ) );
    inv_1 \I6/U1664/U33/U30/Uinv  ( .x(\I6/U1664/U33/Z ), .a(\I6/U1664/y[0] )
         );
    aoi222_1 \I6/U1664/U30/U30/U1  ( .x(\I6/U1664/y[1] ), .a(\I6/U1664/x[3] ), 
        .b(\I6/U1664/x[2] ), .c(\I6/U1664/x[3] ), .d(\I6/U1664/U30/Z ), .e(
        \I6/U1664/x[2] ), .f(\I6/U1664/U30/Z ) );
    inv_1 \I6/U1664/U30/U30/Uinv  ( .x(\I6/U1664/U30/Z ), .a(\I6/U1664/y[1] )
         );
    aoi222_1 \I6/U1664/U31/U30/U1  ( .x(\I6/U1664/x[1] ), .a(\I6/ncd[3] ), .b(
        \I6/ncd[2] ), .c(\I6/ncd[3] ), .d(\I6/U1664/U31/Z ), .e(\I6/ncd[2] ), 
        .f(\I6/U1664/U31/Z ) );
    inv_1 \I6/U1664/U31/U30/Uinv  ( .x(\I6/U1664/U31/Z ), .a(\I6/U1664/x[1] )
         );
    aoi222_1 \I6/U1664/U37/U30/U1  ( .x(\I6/localcd ), .a(\I6/U1664/y[0] ), 
        .b(\I6/U1664/y[1] ), .c(\I6/U1664/y[0] ), .d(\I6/U1664/U37/Z ), .e(
        \I6/U1664/y[1] ), .f(\I6/U1664/U37/Z ) );
    inv_1 \I6/U1664/U37/U30/Uinv  ( .x(\I6/U1664/U37/Z ), .a(\I6/localcd ) );
    nor3_1 \I6/U1669/Unr  ( .x(\I6/U1669/nr ), .a(\I6/ctrlack_internal ), .b(
        n13), .c(\I6/drivel ) );
    nand3_1 \I6/U1669/Und  ( .x(\I6/U1669/nd ), .a(\I6/ctrlack_internal ), .b(
        \I6/driveh ), .c(\I6/drivel ) );
    oa21_1 \I6/U1669/U1  ( .x(\I6/U1669/n2 ), .a(\I6/U1669/n2 ), .b(
        \I6/U1669/nr ), .c(\I6/U1669/nd ) );
    inv_2 \I6/U1669/U3  ( .x(net149), .a(\I6/U1669/n2 ) );
    buf_2 \U1667/U1653  ( .x(\U1667/latch ), .a(net167) );
    nor2_1 \U1667/U264/U5  ( .x(\U1667/nlocalcd ), .a(reset), .b(
        \U1667/localcd ) );
    nor2_1 \U1667/U1659_0_/U5  ( .x(\U1667/ncd[0] ), .a(rd[0]), .b(rd[32]) );
    nor2_1 \U1667/U1659_1_/U5  ( .x(\U1667/ncd[1] ), .a(rd[1]), .b(rd[33]) );
    nor2_1 \U1667/U1659_2_/U5  ( .x(\U1667/ncd[2] ), .a(rd[2]), .b(rd[34]) );
    nor2_1 \U1667/U1659_3_/U5  ( .x(\U1667/ncd[3] ), .a(rd[3]), .b(rd[35]) );
    nor2_1 \U1667/U1659_4_/U5  ( .x(\U1667/ncd[4] ), .a(rd[4]), .b(rd[36]) );
    nor2_1 \U1667/U1659_5_/U5  ( .x(\U1667/ncd[5] ), .a(rd[5]), .b(rd[37]) );
    nor2_1 \U1667/U1659_6_/U5  ( .x(\U1667/ncd[6] ), .a(rd[6]), .b(rd[38]) );
    nor2_1 \U1667/U1659_7_/U5  ( .x(\U1667/ncd[7] ), .a(rd[7]), .b(rd[39]) );
    nor2_1 \U1667/U3/U5  ( .x(\U1667/ctrlack_internal ), .a(\U1667/acb ), .b(
        \U1667/ba ) );
    buf_2 \U1667/U1665/U7  ( .x(\U1667/driveh ), .a(read_lhw) );
    buf_2 \U1667/U1666/U7  ( .x(\U1667/drivel ), .a(read_lhw) );
    ao23_1 \U1667/U1658_0_/U21/U1/U1  ( .x(rd[0]), .a(n11), .b(rd[0]), .c(
        \U1667/drivel ), .d(cbl[0]), .e(n10) );
    ao23_1 \U1667/U1658_1_/U21/U1/U1  ( .x(rd[1]), .a(n11), .b(rd[1]), .c(
        \U1667/driveh ), .d(cbl[1]), .e(n10) );
    ao23_1 \U1667/U1658_2_/U21/U1/U1  ( .x(rd[2]), .a(\U1667/driveh ), .b(rd
        [2]), .c(n11), .d(cbl[2]), .e(n10) );
    ao23_1 \U1667/U1658_3_/U21/U1/U1  ( .x(rd[3]), .a(n11), .b(rd[3]), .c(
        \U1667/driveh ), .d(cbl[3]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_4_/U21/U1/U1  ( .x(rd[4]), .a(\U1667/drivel ), .b(rd
        [4]), .c(n11), .d(cbl[4]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_5_/U21/U1/U1  ( .x(rd[5]), .a(\U1667/drivel ), .b(rd
        [5]), .c(n11), .d(cbl[5]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_6_/U21/U1/U1  ( .x(rd[6]), .a(\U1667/driveh ), .b(rd
        [6]), .c(\U1667/drivel ), .d(cbl[6]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_7_/U21/U1/U1  ( .x(rd[7]), .a(\U1667/driveh ), .b(rd
        [7]), .c(\U1667/driveh ), .d(cbl[7]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_0_/U21/U1/U1  ( .x(rd[32]), .a(\U1667/drivel ), .b(rd
        [32]), .c(n11), .d(cbh[0]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_1_/U21/U1/U1  ( .x(rd[33]), .a(\U1667/driveh ), .b(rd
        [33]), .c(\U1667/drivel ), .d(cbh[1]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_2_/U21/U1/U1  ( .x(rd[34]), .a(\U1667/drivel ), .b(rd
        [34]), .c(\U1667/drivel ), .d(cbh[2]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_3_/U21/U1/U1  ( .x(rd[35]), .a(\U1667/driveh ), .b(rd
        [35]), .c(\U1667/driveh ), .d(cbh[3]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_4_/U21/U1/U1  ( .x(rd[36]), .a(\U1667/drivel ), .b(rd
        [36]), .c(\U1667/driveh ), .d(cbh[4]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_5_/U21/U1/U1  ( .x(rd[37]), .a(\U1667/driveh ), .b(rd
        [37]), .c(n11), .d(cbh[5]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_6_/U21/U1/U1  ( .x(rd[38]), .a(n11), .b(rd[38]), .c(
        \U1667/drivel ), .d(cbh[6]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_7_/U21/U1/U1  ( .x(rd[39]), .a(n11), .b(rd[39]), .c(
        n11), .d(cbh[7]), .e(\U1667/latch ) );
    aoai211_1 \U1667/U4/U28/U1/U1  ( .x(\U1667/U4/U28/U1/clr ), .a(read_lhw), 
        .b(\U1667/acb ), .c(\U1667/nlocalcd ), .d(net167) );
    nand3_1 \U1667/U4/U28/U1/U2  ( .x(\U1667/U4/U28/U1/set ), .a(
        \U1667/nlocalcd ), .b(read_lhw), .c(\U1667/acb ) );
    nand2_2 \U1667/U4/U28/U1/U3  ( .x(net167), .a(\U1667/U4/U28/U1/clr ), .b(
        \U1667/U4/U28/U1/set ) );
    oai21_1 \U1667/U1/U30/U1/U1  ( .x(\U1667/acb ), .a(\U1667/U1/Z ), .b(
        \U1667/ba ), .c(read_lhw) );
    inv_1 \U1667/U1/U30/U1/U2  ( .x(\U1667/U1/Z ), .a(\U1667/acb ) );
    ao222_1 \U1667/U5/U18/U1/U1  ( .x(\U1667/ba ), .a(\U1667/latch ), .b(n14), 
        .c(\U1667/latch ), .d(\U1667/ba ), .e(n14), .f(\U1667/ba ) );
    aoi222_1 \U1667/U1664/U28/U30/U1  ( .x(\U1667/U1664/x[3] ), .a(
        \U1667/ncd[7] ), .b(\U1667/ncd[6] ), .c(\U1667/ncd[7] ), .d(
        \U1667/U1664/U28/Z ), .e(\U1667/ncd[6] ), .f(\U1667/U1664/U28/Z ) );
    inv_1 \U1667/U1664/U28/U30/Uinv  ( .x(\U1667/U1664/U28/Z ), .a(
        \U1667/U1664/x[3] ) );
    aoi222_1 \U1667/U1664/U32/U30/U1  ( .x(\U1667/U1664/x[0] ), .a(
        \U1667/ncd[1] ), .b(\U1667/ncd[0] ), .c(\U1667/ncd[1] ), .d(
        \U1667/U1664/U32/Z ), .e(\U1667/ncd[0] ), .f(\U1667/U1664/U32/Z ) );
    inv_1 \U1667/U1664/U32/U30/Uinv  ( .x(\U1667/U1664/U32/Z ), .a(
        \U1667/U1664/x[0] ) );
    aoi222_1 \U1667/U1664/U29/U30/U1  ( .x(\U1667/U1664/x[2] ), .a(
        \U1667/ncd[5] ), .b(\U1667/ncd[4] ), .c(\U1667/ncd[5] ), .d(
        \U1667/U1664/U29/Z ), .e(\U1667/ncd[4] ), .f(\U1667/U1664/U29/Z ) );
    inv_1 \U1667/U1664/U29/U30/Uinv  ( .x(\U1667/U1664/U29/Z ), .a(
        \U1667/U1664/x[2] ) );
    aoi222_1 \U1667/U1664/U33/U30/U1  ( .x(\U1667/U1664/y[0] ), .a(
        \U1667/U1664/x[1] ), .b(\U1667/U1664/x[0] ), .c(\U1667/U1664/x[1] ), 
        .d(\U1667/U1664/U33/Z ), .e(\U1667/U1664/x[0] ), .f(
        \U1667/U1664/U33/Z ) );
    inv_1 \U1667/U1664/U33/U30/Uinv  ( .x(\U1667/U1664/U33/Z ), .a(
        \U1667/U1664/y[0] ) );
    aoi222_1 \U1667/U1664/U30/U30/U1  ( .x(\U1667/U1664/y[1] ), .a(
        \U1667/U1664/x[3] ), .b(\U1667/U1664/x[2] ), .c(\U1667/U1664/x[3] ), 
        .d(\U1667/U1664/U30/Z ), .e(\U1667/U1664/x[2] ), .f(
        \U1667/U1664/U30/Z ) );
    inv_1 \U1667/U1664/U30/U30/Uinv  ( .x(\U1667/U1664/U30/Z ), .a(
        \U1667/U1664/y[1] ) );
    aoi222_1 \U1667/U1664/U31/U30/U1  ( .x(\U1667/U1664/x[1] ), .a(
        \U1667/ncd[3] ), .b(\U1667/ncd[2] ), .c(\U1667/ncd[3] ), .d(
        \U1667/U1664/U31/Z ), .e(\U1667/ncd[2] ), .f(\U1667/U1664/U31/Z ) );
    inv_1 \U1667/U1664/U31/U30/Uinv  ( .x(\U1667/U1664/U31/Z ), .a(
        \U1667/U1664/x[1] ) );
    aoi222_1 \U1667/U1664/U37/U30/U1  ( .x(\U1667/localcd ), .a(
        \U1667/U1664/y[0] ), .b(\U1667/U1664/y[1] ), .c(\U1667/U1664/y[0] ), 
        .d(\U1667/U1664/U37/Z ), .e(\U1667/U1664/y[1] ), .f(
        \U1667/U1664/U37/Z ) );
    inv_1 \U1667/U1664/U37/U30/Uinv  ( .x(\U1667/U1664/U37/Z ), .a(
        \U1667/localcd ) );
    nor3_1 \U1667/U1669/Unr  ( .x(\U1667/U1669/nr ), .a(
        \U1667/ctrlack_internal ), .b(n11), .c(\U1667/drivel ) );
    nand3_1 \U1667/U1669/Und  ( .x(\U1667/U1669/nd ), .a(
        \U1667/ctrlack_internal ), .b(\U1667/driveh ), .c(\U1667/drivel ) );
    oa21_1 \U1667/U1669/U1  ( .x(\U1667/U1669/n2 ), .a(\U1667/U1669/n2 ), .b(
        \U1667/U1669/nr ), .c(\U1667/U1669/nd ) );
    inv_2 \U1667/U1669/U3  ( .x(net193), .a(\U1667/U1669/n2 ) );
    buf_2 \U1650/U1653  ( .x(\U1650/latch ), .a(net172) );
    nor2_1 \U1650/U264/U5  ( .x(\U1650/nlocalcd ), .a(reset), .b(
        \U1650/localcd ) );
    nor2_1 \U1650/U1659_0_/U5  ( .x(\U1650/ncd[0] ), .a(\U1650/ol[0] ), .b(
        \U1650/oh[0] ) );
    nor2_1 \U1650/U1659_1_/U5  ( .x(\U1650/ncd[1] ), .a(\U1650/ol[1] ), .b(
        \U1650/oh[1] ) );
    nor2_1 \U1650/U1659_2_/U5  ( .x(\U1650/ncd[2] ), .a(\U1650/ol[2] ), .b(
        \U1650/oh[2] ) );
    nor2_1 \U1650/U1659_3_/U5  ( .x(\U1650/ncd[3] ), .a(\U1650/ol[3] ), .b(
        \U1650/oh[3] ) );
    nor2_1 \U1650/U1659_4_/U5  ( .x(\U1650/ncd[4] ), .a(\U1650/ol[4] ), .b(
        \U1650/oh[4] ) );
    nor2_1 \U1650/U1659_5_/U5  ( .x(\U1650/ncd[5] ), .a(\col_l[0] ), .b(
        \col_h[0] ) );
    nor2_1 \U1650/U1659_6_/U5  ( .x(\U1650/ncd[6] ), .a(\col_l[1] ), .b(
        \col_h[1] ) );
    nor2_1 \U1650/U1659_7_/U5  ( .x(\U1650/ncd[7] ), .a(\col_l[2] ), .b(
        \col_h[2] ) );
    nor2_1 \U1650/U3/U5  ( .x(\U1650/ctrlack_internal ), .a(\U1650/acb ), .b(
        \U1650/ba ) );
    buf_2 \U1650/U1665/U7  ( .x(\U1650/driveh ), .a(start_receiving) );
    buf_2 \U1650/U1666/U7  ( .x(\U1650/drivel ), .a(start_receiving) );
    ao23_1 \U1650/U1658_0_/U21/U1/U1  ( .x(\U1650/ol[0] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[0] ), .c(\U1650/drivel ), .d(cbl[0]), .e(n7) );
    ao23_1 \U1650/U1658_1_/U21/U1/U1  ( .x(\U1650/ol[1] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[1] ), .c(\U1650/drivel ), .d(cbl[1]), .e(n7) );
    ao23_1 \U1650/U1658_2_/U21/U1/U1  ( .x(\U1650/ol[2] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[2] ), .c(\U1650/drivel ), .d(cbl[2]), .e(n7) );
    ao23_1 \U1650/U1658_3_/U21/U1/U1  ( .x(\U1650/ol[3] ), .a(n9), .b(
        \U1650/ol[3] ), .c(\U1650/drivel ), .d(cbl[3]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1658_4_/U21/U1/U1  ( .x(\U1650/ol[4] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[4] ), .c(\U1650/drivel ), .d(cbl[4]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1658_5_/U21/U1/U1  ( .x(\col_l[0] ), .a(\U1650/drivel ), 
        .b(\col_l[0] ), .c(\U1650/drivel ), .d(cbl[5]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1658_6_/U21/U1/U1  ( .x(\col_l[1] ), .a(n9), .b(\col_l[1] ), 
        .c(\U1650/drivel ), .d(cbl[6]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1658_7_/U21/U1/U1  ( .x(\col_l[2] ), .a(n9), .b(\col_l[2] ), 
        .c(\U1650/drivel ), .d(cbl[7]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_0_/U21/U1/U1  ( .x(\U1650/oh[0] ), .a(\U1650/driveh ), 
        .b(\U1650/oh[0] ), .c(\U1650/driveh ), .d(cbh[0]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1651_1_/U21/U1/U1  ( .x(\U1650/oh[1] ), .a(\U1650/driveh ), 
        .b(\U1650/oh[1] ), .c(\U1650/driveh ), .d(cbh[1]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1651_2_/U21/U1/U1  ( .x(\U1650/oh[2] ), .a(\U1650/driveh ), 
        .b(\U1650/oh[2] ), .c(\U1650/driveh ), .d(cbh[2]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1651_3_/U21/U1/U1  ( .x(\U1650/oh[3] ), .a(n8), .b(
        \U1650/oh[3] ), .c(\U1650/driveh ), .d(cbh[3]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_4_/U21/U1/U1  ( .x(\U1650/oh[4] ), .a(n8), .b(
        \U1650/oh[4] ), .c(\U1650/driveh ), .d(cbh[4]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_5_/U21/U1/U1  ( .x(\col_h[0] ), .a(\U1650/driveh ), 
        .b(\col_h[0] ), .c(\U1650/driveh ), .d(cbh[5]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_6_/U21/U1/U1  ( .x(\col_h[1] ), .a(n8), .b(\col_h[1] ), 
        .c(\U1650/driveh ), .d(cbh[6]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_7_/U21/U1/U1  ( .x(\col_h[2] ), .a(\U1650/driveh ), 
        .b(\col_h[2] ), .c(\U1650/driveh ), .d(cbh[7]), .e(\U1650/latch ) );
    aoai211_1 \U1650/U4/U28/U1/U1  ( .x(\U1650/U4/U28/U1/clr ), .a(
        start_receiving), .b(\U1650/acb ), .c(\U1650/nlocalcd ), .d(net172) );
    nand3_1 \U1650/U4/U28/U1/U2  ( .x(\U1650/U4/U28/U1/set ), .a(
        \U1650/nlocalcd ), .b(start_receiving), .c(\U1650/acb ) );
    nand2_2 \U1650/U4/U28/U1/U3  ( .x(net172), .a(\U1650/U4/U28/U1/clr ), .b(
        \U1650/U4/U28/U1/set ) );
    oai21_1 \U1650/U1/U30/U1/U1  ( .x(\U1650/acb ), .a(\U1650/U1/Z ), .b(
        \U1650/ba ), .c(start_receiving) );
    inv_1 \U1650/U1/U30/U1/U2  ( .x(\U1650/U1/Z ), .a(\U1650/acb ) );
    ao222_1 \U1650/U5/U18/U1/U1  ( .x(\U1650/ba ), .a(\U1650/latch ), .b(n14), 
        .c(\U1650/latch ), .d(\U1650/ba ), .e(n14), .f(\U1650/ba ) );
    aoi222_1 \U1650/U1664/U28/U30/U1  ( .x(\U1650/U1664/x[3] ), .a(
        \U1650/ncd[7] ), .b(\U1650/ncd[6] ), .c(\U1650/ncd[7] ), .d(
        \U1650/U1664/U28/Z ), .e(\U1650/ncd[6] ), .f(\U1650/U1664/U28/Z ) );
    inv_1 \U1650/U1664/U28/U30/Uinv  ( .x(\U1650/U1664/U28/Z ), .a(
        \U1650/U1664/x[3] ) );
    aoi222_1 \U1650/U1664/U32/U30/U1  ( .x(\U1650/U1664/x[0] ), .a(
        \U1650/ncd[1] ), .b(\U1650/ncd[0] ), .c(\U1650/ncd[1] ), .d(
        \U1650/U1664/U32/Z ), .e(\U1650/ncd[0] ), .f(\U1650/U1664/U32/Z ) );
    inv_1 \U1650/U1664/U32/U30/Uinv  ( .x(\U1650/U1664/U32/Z ), .a(
        \U1650/U1664/x[0] ) );
    aoi222_1 \U1650/U1664/U29/U30/U1  ( .x(\U1650/U1664/x[2] ), .a(
        \U1650/ncd[5] ), .b(\U1650/ncd[4] ), .c(\U1650/ncd[5] ), .d(
        \U1650/U1664/U29/Z ), .e(\U1650/ncd[4] ), .f(\U1650/U1664/U29/Z ) );
    inv_1 \U1650/U1664/U29/U30/Uinv  ( .x(\U1650/U1664/U29/Z ), .a(
        \U1650/U1664/x[2] ) );
    aoi222_1 \U1650/U1664/U33/U30/U1  ( .x(\U1650/U1664/y[0] ), .a(
        \U1650/U1664/x[1] ), .b(\U1650/U1664/x[0] ), .c(\U1650/U1664/x[1] ), 
        .d(\U1650/U1664/U33/Z ), .e(\U1650/U1664/x[0] ), .f(
        \U1650/U1664/U33/Z ) );
    inv_1 \U1650/U1664/U33/U30/Uinv  ( .x(\U1650/U1664/U33/Z ), .a(
        \U1650/U1664/y[0] ) );
    aoi222_1 \U1650/U1664/U30/U30/U1  ( .x(\U1650/U1664/y[1] ), .a(
        \U1650/U1664/x[3] ), .b(\U1650/U1664/x[2] ), .c(\U1650/U1664/x[3] ), 
        .d(\U1650/U1664/U30/Z ), .e(\U1650/U1664/x[2] ), .f(
        \U1650/U1664/U30/Z ) );
    inv_1 \U1650/U1664/U30/U30/Uinv  ( .x(\U1650/U1664/U30/Z ), .a(
        \U1650/U1664/y[1] ) );
    aoi222_1 \U1650/U1664/U31/U30/U1  ( .x(\U1650/U1664/x[1] ), .a(
        \U1650/ncd[3] ), .b(\U1650/ncd[2] ), .c(\U1650/ncd[3] ), .d(
        \U1650/U1664/U31/Z ), .e(\U1650/ncd[2] ), .f(\U1650/U1664/U31/Z ) );
    inv_1 \U1650/U1664/U31/U30/Uinv  ( .x(\U1650/U1664/U31/Z ), .a(
        \U1650/U1664/x[1] ) );
    aoi222_1 \U1650/U1664/U37/U30/U1  ( .x(\U1650/localcd ), .a(
        \U1650/U1664/y[0] ), .b(\U1650/U1664/y[1] ), .c(\U1650/U1664/y[0] ), 
        .d(\U1650/U1664/U37/Z ), .e(\U1650/U1664/y[1] ), .f(
        \U1650/U1664/U37/Z ) );
    inv_1 \U1650/U1664/U37/U30/Uinv  ( .x(\U1650/U1664/U37/Z ), .a(
        \U1650/localcd ) );
    nor3_1 \U1650/U1669/Unr  ( .x(\U1650/U1669/nr ), .a(
        \U1650/ctrlack_internal ), .b(\U1650/drivel ), .c(\U1650/driveh ) );
    nand3_1 \U1650/U1669/Und  ( .x(\U1650/U1669/nd ), .a(
        \U1650/ctrlack_internal ), .b(\U1650/drivel ), .c(\U1650/driveh ) );
    oa21_1 \U1650/U1669/U1  ( .x(\U1650/U1669/n2 ), .a(\U1650/U1669/n2 ), .b(
        \U1650/U1669/nr ), .c(\U1650/U1669/nd ) );
    inv_2 \U1650/U1669/U3  ( .x(net139), .a(\U1650/U1669/n2 ) );
    buf_2 \U1666/U1653  ( .x(\U1666/latch ), .a(net169) );
    nor2_1 \U1666/U264/U5  ( .x(\U1666/nlocalcd ), .a(reset), .b(
        \U1666/localcd ) );
    nor2_1 \U1666/U1659_0_/U5  ( .x(\U1666/ncd[0] ), .a(rd[24]), .b(rd[56]) );
    nor2_1 \U1666/U1659_1_/U5  ( .x(\U1666/ncd[1] ), .a(rd[25]), .b(rd[57]) );
    nor2_1 \U1666/U1659_2_/U5  ( .x(\U1666/ncd[2] ), .a(rd[26]), .b(rd[58]) );
    nor2_1 \U1666/U1659_3_/U5  ( .x(\U1666/ncd[3] ), .a(rd[27]), .b(rd[59]) );
    nor2_1 \U1666/U1659_4_/U5  ( .x(\U1666/ncd[4] ), .a(rd[28]), .b(rd[60]) );
    nor2_1 \U1666/U1659_5_/U5  ( .x(\U1666/ncd[5] ), .a(rd[29]), .b(rd[61]) );
    nor2_1 \U1666/U1659_6_/U5  ( .x(\U1666/ncd[6] ), .a(rd[30]), .b(rd[62]) );
    nor2_1 \U1666/U1659_7_/U5  ( .x(\U1666/ncd[7] ), .a(rd[31]), .b(rd[63]) );
    nor2_1 \U1666/U3/U5  ( .x(\U1666/ctrlack_internal ), .a(\U1666/acb ), .b(
        \U1666/ba ) );
    buf_2 \U1666/U1665/U7  ( .x(\U1666/driveh ), .a(read) );
    buf_2 \U1666/U1666/U7  ( .x(\U1666/drivel ), .a(read) );
    ao23_1 \U1666/U1658_0_/U21/U1/U1  ( .x(rd[24]), .a(n6), .b(rd[24]), .c(
        \U1666/drivel ), .d(cbl[0]), .e(n5) );
    ao23_1 \U1666/U1658_1_/U21/U1/U1  ( .x(rd[25]), .a(n6), .b(rd[25]), .c(
        \U1666/driveh ), .d(cbl[1]), .e(n5) );
    ao23_1 \U1666/U1658_2_/U21/U1/U1  ( .x(rd[26]), .a(\U1666/driveh ), .b(rd
        [26]), .c(n6), .d(cbl[2]), .e(n5) );
    ao23_1 \U1666/U1658_3_/U21/U1/U1  ( .x(rd[27]), .a(n6), .b(rd[27]), .c(
        \U1666/driveh ), .d(cbl[3]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_4_/U21/U1/U1  ( .x(rd[28]), .a(\U1666/drivel ), .b(rd
        [28]), .c(n6), .d(cbl[4]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_5_/U21/U1/U1  ( .x(rd[29]), .a(\U1666/drivel ), .b(rd
        [29]), .c(n6), .d(cbl[5]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_6_/U21/U1/U1  ( .x(rd[30]), .a(\U1666/driveh ), .b(rd
        [30]), .c(\U1666/drivel ), .d(cbl[6]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_7_/U21/U1/U1  ( .x(rd[31]), .a(\U1666/driveh ), .b(rd
        [31]), .c(\U1666/driveh ), .d(cbl[7]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_0_/U21/U1/U1  ( .x(rd[56]), .a(\U1666/drivel ), .b(rd
        [56]), .c(n6), .d(cbh[0]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_1_/U21/U1/U1  ( .x(rd[57]), .a(\U1666/driveh ), .b(rd
        [57]), .c(\U1666/drivel ), .d(cbh[1]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_2_/U21/U1/U1  ( .x(rd[58]), .a(\U1666/drivel ), .b(rd
        [58]), .c(\U1666/drivel ), .d(cbh[2]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_3_/U21/U1/U1  ( .x(rd[59]), .a(\U1666/driveh ), .b(rd
        [59]), .c(\U1666/driveh ), .d(cbh[3]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_4_/U21/U1/U1  ( .x(rd[60]), .a(\U1666/drivel ), .b(rd
        [60]), .c(\U1666/driveh ), .d(cbh[4]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_5_/U21/U1/U1  ( .x(rd[61]), .a(\U1666/driveh ), .b(rd
        [61]), .c(n6), .d(cbh[5]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_6_/U21/U1/U1  ( .x(rd[62]), .a(n6), .b(rd[62]), .c(
        \U1666/drivel ), .d(cbh[6]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_7_/U21/U1/U1  ( .x(rd[63]), .a(n6), .b(rd[63]), .c(n6), 
        .d(cbh[7]), .e(\U1666/latch ) );
    aoai211_1 \U1666/U4/U28/U1/U1  ( .x(\U1666/U4/U28/U1/clr ), .a(read), .b(
        \U1666/acb ), .c(\U1666/nlocalcd ), .d(net169) );
    nand3_1 \U1666/U4/U28/U1/U2  ( .x(\U1666/U4/U28/U1/set ), .a(
        \U1666/nlocalcd ), .b(read), .c(\U1666/acb ) );
    nand2_2 \U1666/U4/U28/U1/U3  ( .x(net169), .a(\U1666/U4/U28/U1/clr ), .b(
        \U1666/U4/U28/U1/set ) );
    oai21_1 \U1666/U1/U30/U1/U1  ( .x(\U1666/acb ), .a(\U1666/U1/Z ), .b(
        \U1666/ba ), .c(read) );
    inv_1 \U1666/U1/U30/U1/U2  ( .x(\U1666/U1/Z ), .a(\U1666/acb ) );
    ao222_1 \U1666/U5/U18/U1/U1  ( .x(\U1666/ba ), .a(\U1666/latch ), .b(n14), 
        .c(\U1666/latch ), .d(\U1666/ba ), .e(n14), .f(\U1666/ba ) );
    aoi222_1 \U1666/U1664/U28/U30/U1  ( .x(\U1666/U1664/x[3] ), .a(
        \U1666/ncd[7] ), .b(\U1666/ncd[6] ), .c(\U1666/ncd[7] ), .d(
        \U1666/U1664/U28/Z ), .e(\U1666/ncd[6] ), .f(\U1666/U1664/U28/Z ) );
    inv_1 \U1666/U1664/U28/U30/Uinv  ( .x(\U1666/U1664/U28/Z ), .a(
        \U1666/U1664/x[3] ) );
    aoi222_1 \U1666/U1664/U32/U30/U1  ( .x(\U1666/U1664/x[0] ), .a(
        \U1666/ncd[1] ), .b(\U1666/ncd[0] ), .c(\U1666/ncd[1] ), .d(
        \U1666/U1664/U32/Z ), .e(\U1666/ncd[0] ), .f(\U1666/U1664/U32/Z ) );
    inv_1 \U1666/U1664/U32/U30/Uinv  ( .x(\U1666/U1664/U32/Z ), .a(
        \U1666/U1664/x[0] ) );
    aoi222_1 \U1666/U1664/U29/U30/U1  ( .x(\U1666/U1664/x[2] ), .a(
        \U1666/ncd[5] ), .b(\U1666/ncd[4] ), .c(\U1666/ncd[5] ), .d(
        \U1666/U1664/U29/Z ), .e(\U1666/ncd[4] ), .f(\U1666/U1664/U29/Z ) );
    inv_1 \U1666/U1664/U29/U30/Uinv  ( .x(\U1666/U1664/U29/Z ), .a(
        \U1666/U1664/x[2] ) );
    aoi222_1 \U1666/U1664/U33/U30/U1  ( .x(\U1666/U1664/y[0] ), .a(
        \U1666/U1664/x[1] ), .b(\U1666/U1664/x[0] ), .c(\U1666/U1664/x[1] ), 
        .d(\U1666/U1664/U33/Z ), .e(\U1666/U1664/x[0] ), .f(
        \U1666/U1664/U33/Z ) );
    inv_1 \U1666/U1664/U33/U30/Uinv  ( .x(\U1666/U1664/U33/Z ), .a(
        \U1666/U1664/y[0] ) );
    aoi222_1 \U1666/U1664/U30/U30/U1  ( .x(\U1666/U1664/y[1] ), .a(
        \U1666/U1664/x[3] ), .b(\U1666/U1664/x[2] ), .c(\U1666/U1664/x[3] ), 
        .d(\U1666/U1664/U30/Z ), .e(\U1666/U1664/x[2] ), .f(
        \U1666/U1664/U30/Z ) );
    inv_1 \U1666/U1664/U30/U30/Uinv  ( .x(\U1666/U1664/U30/Z ), .a(
        \U1666/U1664/y[1] ) );
    aoi222_1 \U1666/U1664/U31/U30/U1  ( .x(\U1666/U1664/x[1] ), .a(
        \U1666/ncd[3] ), .b(\U1666/ncd[2] ), .c(\U1666/ncd[3] ), .d(
        \U1666/U1664/U31/Z ), .e(\U1666/ncd[2] ), .f(\U1666/U1664/U31/Z ) );
    inv_1 \U1666/U1664/U31/U30/Uinv  ( .x(\U1666/U1664/U31/Z ), .a(
        \U1666/U1664/x[1] ) );
    aoi222_1 \U1666/U1664/U37/U30/U1  ( .x(\U1666/localcd ), .a(
        \U1666/U1664/y[0] ), .b(\U1666/U1664/y[1] ), .c(\U1666/U1664/y[0] ), 
        .d(\U1666/U1664/U37/Z ), .e(\U1666/U1664/y[1] ), .f(
        \U1666/U1664/U37/Z ) );
    inv_1 \U1666/U1664/U37/U30/Uinv  ( .x(\U1666/U1664/U37/Z ), .a(
        \U1666/localcd ) );
    nor3_1 \U1666/U1669/Unr  ( .x(\U1666/U1669/nr ), .a(
        \U1666/ctrlack_internal ), .b(n6), .c(\U1666/drivel ) );
    nand3_1 \U1666/U1669/Und  ( .x(\U1666/U1669/nd ), .a(
        \U1666/ctrlack_internal ), .b(\U1666/driveh ), .c(\U1666/drivel ) );
    oa21_1 \U1666/U1669/U1  ( .x(\U1666/U1669/n2 ), .a(\U1666/U1669/n2 ), .b(
        \U1666/U1669/nr ), .c(\U1666/U1669/nd ) );
    inv_2 \U1666/U1669/U3  ( .x(net94), .a(\U1666/U1669/n2 ) );
    buf_2 \I1/U1653  ( .x(\I1/latch ), .a(net166) );
    nor2_1 \I1/U264/U5  ( .x(\I1/nlocalcd ), .a(reset), .b(\I1/localcd ) );
    nor2_1 \I1/U1659_0_/U5  ( .x(\I1/ncd[0] ), .a(rd[8]), .b(rd[40]) );
    nor2_1 \I1/U1659_1_/U5  ( .x(\I1/ncd[1] ), .a(rd[9]), .b(rd[41]) );
    nor2_1 \I1/U1659_2_/U5  ( .x(\I1/ncd[2] ), .a(rd[10]), .b(rd[42]) );
    nor2_1 \I1/U1659_3_/U5  ( .x(\I1/ncd[3] ), .a(rd[11]), .b(rd[43]) );
    nor2_1 \I1/U1659_4_/U5  ( .x(\I1/ncd[4] ), .a(rd[12]), .b(rd[44]) );
    nor2_1 \I1/U1659_5_/U5  ( .x(\I1/ncd[5] ), .a(rd[13]), .b(rd[45]) );
    nor2_1 \I1/U1659_6_/U5  ( .x(\I1/ncd[6] ), .a(rd[14]), .b(rd[46]) );
    nor2_1 \I1/U1659_7_/U5  ( .x(\I1/ncd[7] ), .a(rd[15]), .b(rd[47]) );
    nor2_1 \I1/U3/U5  ( .x(\I1/ctrlack_internal ), .a(\I1/acb ), .b(\I1/ba )
         );
    buf_2 \I1/U1665/U7  ( .x(\I1/driveh ), .a(net103) );
    buf_2 \I1/U1666/U7  ( .x(\I1/drivel ), .a(net103) );
    ao23_1 \I1/U1658_0_/U21/U1/U1  ( .x(rd[8]), .a(n4), .b(rd[8]), .c(
        \I1/drivel ), .d(cbl[0]), .e(n3) );
    ao23_1 \I1/U1658_1_/U21/U1/U1  ( .x(rd[9]), .a(n4), .b(rd[9]), .c(
        \I1/driveh ), .d(cbl[1]), .e(n3) );
    ao23_1 \I1/U1658_2_/U21/U1/U1  ( .x(rd[10]), .a(\I1/driveh ), .b(rd[10]), 
        .c(n4), .d(cbl[2]), .e(n3) );
    ao23_1 \I1/U1658_3_/U21/U1/U1  ( .x(rd[11]), .a(n4), .b(rd[11]), .c(
        \I1/driveh ), .d(cbl[3]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_4_/U21/U1/U1  ( .x(rd[12]), .a(\I1/drivel ), .b(rd[12]), 
        .c(n4), .d(cbl[4]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_5_/U21/U1/U1  ( .x(rd[13]), .a(\I1/drivel ), .b(rd[13]), 
        .c(n4), .d(cbl[5]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_6_/U21/U1/U1  ( .x(rd[14]), .a(\I1/driveh ), .b(rd[14]), 
        .c(\I1/drivel ), .d(cbl[6]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_7_/U21/U1/U1  ( .x(rd[15]), .a(\I1/driveh ), .b(rd[15]), 
        .c(\I1/driveh ), .d(cbl[7]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_0_/U21/U1/U1  ( .x(rd[40]), .a(\I1/drivel ), .b(rd[40]), 
        .c(n4), .d(cbh[0]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_1_/U21/U1/U1  ( .x(rd[41]), .a(\I1/driveh ), .b(rd[41]), 
        .c(\I1/drivel ), .d(cbh[1]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_2_/U21/U1/U1  ( .x(rd[42]), .a(\I1/drivel ), .b(rd[42]), 
        .c(\I1/drivel ), .d(cbh[2]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_3_/U21/U1/U1  ( .x(rd[43]), .a(\I1/driveh ), .b(rd[43]), 
        .c(\I1/driveh ), .d(cbh[3]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_4_/U21/U1/U1  ( .x(rd[44]), .a(\I1/drivel ), .b(rd[44]), 
        .c(\I1/driveh ), .d(cbh[4]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_5_/U21/U1/U1  ( .x(rd[45]), .a(\I1/driveh ), .b(rd[45]), 
        .c(n4), .d(cbh[5]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_6_/U21/U1/U1  ( .x(rd[46]), .a(n4), .b(rd[46]), .c(
        \I1/drivel ), .d(cbh[6]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_7_/U21/U1/U1  ( .x(rd[47]), .a(n4), .b(rd[47]), .c(n4), 
        .d(cbh[7]), .e(\I1/latch ) );
    aoai211_1 \I1/U4/U28/U1/U1  ( .x(\I1/U4/U28/U1/clr ), .a(net103), .b(
        \I1/acb ), .c(\I1/nlocalcd ), .d(net166) );
    nand3_1 \I1/U4/U28/U1/U2  ( .x(\I1/U4/U28/U1/set ), .a(\I1/nlocalcd ), .b(
        net103), .c(\I1/acb ) );
    nand2_2 \I1/U4/U28/U1/U3  ( .x(net166), .a(\I1/U4/U28/U1/clr ), .b(
        \I1/U4/U28/U1/set ) );
    oai21_1 \I1/U1/U30/U1/U1  ( .x(\I1/acb ), .a(\I1/U1/Z ), .b(\I1/ba ), .c(
        net103) );
    inv_1 \I1/U1/U30/U1/U2  ( .x(\I1/U1/Z ), .a(\I1/acb ) );
    ao222_1 \I1/U5/U18/U1/U1  ( .x(\I1/ba ), .a(\I1/latch ), .b(n14), .c(
        \I1/latch ), .d(\I1/ba ), .e(n14), .f(\I1/ba ) );
    aoi222_1 \I1/U1664/U28/U30/U1  ( .x(\I1/U1664/x[3] ), .a(\I1/ncd[7] ), .b(
        \I1/ncd[6] ), .c(\I1/ncd[7] ), .d(\I1/U1664/U28/Z ), .e(\I1/ncd[6] ), 
        .f(\I1/U1664/U28/Z ) );
    inv_1 \I1/U1664/U28/U30/Uinv  ( .x(\I1/U1664/U28/Z ), .a(\I1/U1664/x[3] )
         );
    aoi222_1 \I1/U1664/U32/U30/U1  ( .x(\I1/U1664/x[0] ), .a(\I1/ncd[1] ), .b(
        \I1/ncd[0] ), .c(\I1/ncd[1] ), .d(\I1/U1664/U32/Z ), .e(\I1/ncd[0] ), 
        .f(\I1/U1664/U32/Z ) );
    inv_1 \I1/U1664/U32/U30/Uinv  ( .x(\I1/U1664/U32/Z ), .a(\I1/U1664/x[0] )
         );
    aoi222_1 \I1/U1664/U29/U30/U1  ( .x(\I1/U1664/x[2] ), .a(\I1/ncd[5] ), .b(
        \I1/ncd[4] ), .c(\I1/ncd[5] ), .d(\I1/U1664/U29/Z ), .e(\I1/ncd[4] ), 
        .f(\I1/U1664/U29/Z ) );
    inv_1 \I1/U1664/U29/U30/Uinv  ( .x(\I1/U1664/U29/Z ), .a(\I1/U1664/x[2] )
         );
    aoi222_1 \I1/U1664/U33/U30/U1  ( .x(\I1/U1664/y[0] ), .a(\I1/U1664/x[1] ), 
        .b(\I1/U1664/x[0] ), .c(\I1/U1664/x[1] ), .d(\I1/U1664/U33/Z ), .e(
        \I1/U1664/x[0] ), .f(\I1/U1664/U33/Z ) );
    inv_1 \I1/U1664/U33/U30/Uinv  ( .x(\I1/U1664/U33/Z ), .a(\I1/U1664/y[0] )
         );
    aoi222_1 \I1/U1664/U30/U30/U1  ( .x(\I1/U1664/y[1] ), .a(\I1/U1664/x[3] ), 
        .b(\I1/U1664/x[2] ), .c(\I1/U1664/x[3] ), .d(\I1/U1664/U30/Z ), .e(
        \I1/U1664/x[2] ), .f(\I1/U1664/U30/Z ) );
    inv_1 \I1/U1664/U30/U30/Uinv  ( .x(\I1/U1664/U30/Z ), .a(\I1/U1664/y[1] )
         );
    aoi222_1 \I1/U1664/U31/U30/U1  ( .x(\I1/U1664/x[1] ), .a(\I1/ncd[3] ), .b(
        \I1/ncd[2] ), .c(\I1/ncd[3] ), .d(\I1/U1664/U31/Z ), .e(\I1/ncd[2] ), 
        .f(\I1/U1664/U31/Z ) );
    inv_1 \I1/U1664/U31/U30/Uinv  ( .x(\I1/U1664/U31/Z ), .a(\I1/U1664/x[1] )
         );
    aoi222_1 \I1/U1664/U37/U30/U1  ( .x(\I1/localcd ), .a(\I1/U1664/y[0] ), 
        .b(\I1/U1664/y[1] ), .c(\I1/U1664/y[0] ), .d(\I1/U1664/U37/Z ), .e(
        \I1/U1664/y[1] ), .f(\I1/U1664/U37/Z ) );
    inv_1 \I1/U1664/U37/U30/Uinv  ( .x(\I1/U1664/U37/Z ), .a(\I1/localcd ) );
    nor3_1 \I1/U1669/Unr  ( .x(\I1/U1669/nr ), .a(\I1/ctrlack_internal ), .b(
        n4), .c(\I1/drivel ) );
    nand3_1 \I1/U1669/Und  ( .x(\I1/U1669/nd ), .a(\I1/ctrlack_internal ), .b(
        \I1/driveh ), .c(\I1/drivel ) );
    oa21_1 \I1/U1669/U1  ( .x(\I1/U1669/n2 ), .a(\I1/U1669/n2 ), .b(
        \I1/U1669/nr ), .c(\I1/U1669/nd ) );
    inv_2 \I1/U1669/U3  ( .x(read_lhw), .a(\I1/U1669/n2 ) );
    buf_2 \I2/U1653  ( .x(\I2/latch ), .a(net170) );
    nor2_1 \I2/U264/U5  ( .x(\I2/nlocalcd ), .a(reset), .b(\I2/localcd ) );
    nor2_1 \I2/U1659_0_/U5  ( .x(\I2/ncd[0] ), .a(rd[16]), .b(rd[48]) );
    nor2_1 \I2/U1659_1_/U5  ( .x(\I2/ncd[1] ), .a(rd[17]), .b(rd[49]) );
    nor2_1 \I2/U1659_2_/U5  ( .x(\I2/ncd[2] ), .a(rd[18]), .b(rd[50]) );
    nor2_1 \I2/U1659_3_/U5  ( .x(\I2/ncd[3] ), .a(rd[19]), .b(rd[51]) );
    nor2_1 \I2/U1659_4_/U5  ( .x(\I2/ncd[4] ), .a(rd[20]), .b(rd[52]) );
    nor2_1 \I2/U1659_5_/U5  ( .x(\I2/ncd[5] ), .a(rd[21]), .b(rd[53]) );
    nor2_1 \I2/U1659_6_/U5  ( .x(\I2/ncd[6] ), .a(rd[22]), .b(rd[54]) );
    nor2_1 \I2/U1659_7_/U5  ( .x(\I2/ncd[7] ), .a(rd[23]), .b(rd[55]) );
    nor2_1 \I2/U3/U5  ( .x(\I2/ctrlack_internal ), .a(\I2/acb ), .b(\I2/ba )
         );
    buf_2 \I2/U1665/U7  ( .x(\I2/driveh ), .a(net94) );
    buf_2 \I2/U1666/U7  ( .x(\I2/drivel ), .a(net94) );
    ao23_1 \I2/U1658_0_/U21/U1/U1  ( .x(rd[16]), .a(n2), .b(rd[16]), .c(
        \I2/drivel ), .d(cbl[0]), .e(n1) );
    ao23_1 \I2/U1658_1_/U21/U1/U1  ( .x(rd[17]), .a(n2), .b(rd[17]), .c(
        \I2/driveh ), .d(cbl[1]), .e(n1) );
    ao23_1 \I2/U1658_2_/U21/U1/U1  ( .x(rd[18]), .a(\I2/driveh ), .b(rd[18]), 
        .c(n2), .d(cbl[2]), .e(n1) );
    ao23_1 \I2/U1658_3_/U21/U1/U1  ( .x(rd[19]), .a(n2), .b(rd[19]), .c(
        \I2/driveh ), .d(cbl[3]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_4_/U21/U1/U1  ( .x(rd[20]), .a(\I2/drivel ), .b(rd[20]), 
        .c(n2), .d(cbl[4]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_5_/U21/U1/U1  ( .x(rd[21]), .a(\I2/drivel ), .b(rd[21]), 
        .c(n2), .d(cbl[5]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_6_/U21/U1/U1  ( .x(rd[22]), .a(\I2/driveh ), .b(rd[22]), 
        .c(\I2/drivel ), .d(cbl[6]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_7_/U21/U1/U1  ( .x(rd[23]), .a(\I2/driveh ), .b(rd[23]), 
        .c(\I2/driveh ), .d(cbl[7]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_0_/U21/U1/U1  ( .x(rd[48]), .a(\I2/drivel ), .b(rd[48]), 
        .c(n2), .d(cbh[0]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_1_/U21/U1/U1  ( .x(rd[49]), .a(\I2/driveh ), .b(rd[49]), 
        .c(\I2/drivel ), .d(cbh[1]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_2_/U21/U1/U1  ( .x(rd[50]), .a(\I2/drivel ), .b(rd[50]), 
        .c(\I2/drivel ), .d(cbh[2]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_3_/U21/U1/U1  ( .x(rd[51]), .a(\I2/driveh ), .b(rd[51]), 
        .c(\I2/driveh ), .d(cbh[3]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_4_/U21/U1/U1  ( .x(rd[52]), .a(\I2/drivel ), .b(rd[52]), 
        .c(\I2/driveh ), .d(cbh[4]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_5_/U21/U1/U1  ( .x(rd[53]), .a(\I2/driveh ), .b(rd[53]), 
        .c(n2), .d(cbh[5]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_6_/U21/U1/U1  ( .x(rd[54]), .a(n2), .b(rd[54]), .c(
        \I2/drivel ), .d(cbh[6]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_7_/U21/U1/U1  ( .x(rd[55]), .a(n2), .b(rd[55]), .c(n2), 
        .d(cbh[7]), .e(\I2/latch ) );
    aoai211_1 \I2/U4/U28/U1/U1  ( .x(\I2/U4/U28/U1/clr ), .a(net94), .b(
        \I2/acb ), .c(\I2/nlocalcd ), .d(net170) );
    nand3_1 \I2/U4/U28/U1/U2  ( .x(\I2/U4/U28/U1/set ), .a(\I2/nlocalcd ), .b(
        net94), .c(\I2/acb ) );
    nand2_2 \I2/U4/U28/U1/U3  ( .x(net170), .a(\I2/U4/U28/U1/clr ), .b(
        \I2/U4/U28/U1/set ) );
    oai21_1 \I2/U1/U30/U1/U1  ( .x(\I2/acb ), .a(\I2/U1/Z ), .b(\I2/ba ), .c(
        net94) );
    inv_1 \I2/U1/U30/U1/U2  ( .x(\I2/U1/Z ), .a(\I2/acb ) );
    ao222_1 \I2/U5/U18/U1/U1  ( .x(\I2/ba ), .a(\I2/latch ), .b(n14), .c(
        \I2/latch ), .d(\I2/ba ), .e(n14), .f(\I2/ba ) );
    aoi222_1 \I2/U1664/U28/U30/U1  ( .x(\I2/U1664/x[3] ), .a(\I2/ncd[7] ), .b(
        \I2/ncd[6] ), .c(\I2/ncd[7] ), .d(\I2/U1664/U28/Z ), .e(\I2/ncd[6] ), 
        .f(\I2/U1664/U28/Z ) );
    inv_1 \I2/U1664/U28/U30/Uinv  ( .x(\I2/U1664/U28/Z ), .a(\I2/U1664/x[3] )
         );
    aoi222_1 \I2/U1664/U32/U30/U1  ( .x(\I2/U1664/x[0] ), .a(\I2/ncd[1] ), .b(
        \I2/ncd[0] ), .c(\I2/ncd[1] ), .d(\I2/U1664/U32/Z ), .e(\I2/ncd[0] ), 
        .f(\I2/U1664/U32/Z ) );
    inv_1 \I2/U1664/U32/U30/Uinv  ( .x(\I2/U1664/U32/Z ), .a(\I2/U1664/x[0] )
         );
    aoi222_1 \I2/U1664/U29/U30/U1  ( .x(\I2/U1664/x[2] ), .a(\I2/ncd[5] ), .b(
        \I2/ncd[4] ), .c(\I2/ncd[5] ), .d(\I2/U1664/U29/Z ), .e(\I2/ncd[4] ), 
        .f(\I2/U1664/U29/Z ) );
    inv_1 \I2/U1664/U29/U30/Uinv  ( .x(\I2/U1664/U29/Z ), .a(\I2/U1664/x[2] )
         );
    aoi222_1 \I2/U1664/U33/U30/U1  ( .x(\I2/U1664/y[0] ), .a(\I2/U1664/x[1] ), 
        .b(\I2/U1664/x[0] ), .c(\I2/U1664/x[1] ), .d(\I2/U1664/U33/Z ), .e(
        \I2/U1664/x[0] ), .f(\I2/U1664/U33/Z ) );
    inv_1 \I2/U1664/U33/U30/Uinv  ( .x(\I2/U1664/U33/Z ), .a(\I2/U1664/y[0] )
         );
    aoi222_1 \I2/U1664/U30/U30/U1  ( .x(\I2/U1664/y[1] ), .a(\I2/U1664/x[3] ), 
        .b(\I2/U1664/x[2] ), .c(\I2/U1664/x[3] ), .d(\I2/U1664/U30/Z ), .e(
        \I2/U1664/x[2] ), .f(\I2/U1664/U30/Z ) );
    inv_1 \I2/U1664/U30/U30/Uinv  ( .x(\I2/U1664/U30/Z ), .a(\I2/U1664/y[1] )
         );
    aoi222_1 \I2/U1664/U31/U30/U1  ( .x(\I2/U1664/x[1] ), .a(\I2/ncd[3] ), .b(
        \I2/ncd[2] ), .c(\I2/ncd[3] ), .d(\I2/U1664/U31/Z ), .e(\I2/ncd[2] ), 
        .f(\I2/U1664/U31/Z ) );
    inv_1 \I2/U1664/U31/U30/Uinv  ( .x(\I2/U1664/U31/Z ), .a(\I2/U1664/x[1] )
         );
    aoi222_1 \I2/U1664/U37/U30/U1  ( .x(\I2/localcd ), .a(\I2/U1664/y[0] ), 
        .b(\I2/U1664/y[1] ), .c(\I2/U1664/y[0] ), .d(\I2/U1664/U37/Z ), .e(
        \I2/U1664/y[1] ), .f(\I2/U1664/U37/Z ) );
    inv_1 \I2/U1664/U37/U30/Uinv  ( .x(\I2/U1664/U37/Z ), .a(\I2/localcd ) );
    nor3_1 \I2/U1669/Unr  ( .x(\I2/U1669/nr ), .a(\I2/ctrlack_internal ), .b(
        n2), .c(\I2/drivel ) );
    nand3_1 \I2/U1669/Und  ( .x(\I2/U1669/nd ), .a(\I2/ctrlack_internal ), .b(
        \I2/driveh ), .c(\I2/drivel ) );
    oa21_1 \I2/U1669/U1  ( .x(\I2/U1669/n2 ), .a(\I2/U1669/n2 ), .b(
        \I2/U1669/nr ), .c(\I2/U1669/nd ) );
    inv_2 \I2/U1669/U3  ( .x(net103), .a(\I2/U1669/n2 ) );
    buf_1 U1 ( .x(n1), .a(\I2/latch ) );
    buf_2 U2 ( .x(n2), .a(net94) );
    buf_1 U3 ( .x(n3), .a(\I1/latch ) );
    buf_2 U4 ( .x(n4), .a(net103) );
    buf_1 U5 ( .x(n5), .a(\U1666/latch ) );
    buf_2 U6 ( .x(n6), .a(read) );
    buf_1 U7 ( .x(n7), .a(\U1650/latch ) );
    buf_1 U8 ( .x(n8), .a(\U1650/driveh ) );
    buf_1 U9 ( .x(n9), .a(\U1650/drivel ) );
    buf_1 U10 ( .x(n10), .a(\U1667/latch ) );
    buf_2 U11 ( .x(n11), .a(read_lhw) );
    buf_1 U12 ( .x(n12), .a(\I6/latch ) );
    buf_2 U13 ( .x(n13), .a(net139) );
    buf_3 U14 ( .x(n14), .a(bpullcd) );
    buf_3 U15 ( .x(err[0]), .a(n18) );
    buf_3 U16 ( .x(err[1]), .a(n17) );
endmodule


module chain_fr2dr_byte_3 ( nia, oh, ol, i, nReset, noa );
output [7:0] oh;
output [7:0] ol;
input  [4:0] i;
input  nReset, noa;
output nia;
    wire eop, net135, nca, nbReset, ncla, \c[3] , \c[2] , \c[1] , \c[0] , 
        \cl[3] , \cl[2] , \cl[1] , \cl[0] , asel, bsel, asela, bsela, csel, 
        dsel, csela, dsela, esel, fsel, esela, fsela, naa, nda, \a[3] , \a[2] , 
        \a[1] , \a[0] , \d[3] , \d[2] , \d[1] , \d[0] , nba, nea, nfa, \b[3] , 
        \b[2] , \b[1] , \b[0] , \f[3] , \f[2] , \f[1] , \f[0] , \e[3] , \e[2] , 
        \e[1] , \e[0] , \U891/nack , \U891/acka , \U891/naack[0] , 
        \U891/naack[1] , \U891/iay , \U891/ackb , \U891/reset , \U891/neopack , 
        \U891/U1128/nb , \U891/U1128/na , \U891/U1118_0_/nr , 
        \U891/U1118_0_/nd , \U891/U1118_0_/n2 , \U891/U1118_1_/nr , 
        \U891/U1118_1_/nd , \U891/U1118_1_/n2 , \U891/U1118_2_/nr , 
        \U891/U1118_2_/nd , \U891/U1118_2_/n2 , \U891/U1118_3_/nr , 
        \U891/U1118_3_/nd , \U891/U1118_3_/n2 , \U891/U1117_0_/nr , 
        \U891/U1117_0_/nd , \U891/U1117_0_/n2 , \U891/U1117_1_/nr , 
        \U891/U1117_1_/nd , \U891/U1117_1_/n2 , \U891/U1117_2_/nr , 
        \U891/U1117_2_/nd , \U891/U1117_2_/n2 , \U891/U1117_3_/nr , 
        \U891/U1117_3_/nd , \U891/U1117_3_/n2 , \U886/nack , \U886/acka , 
        \U886/ackb , \U886/reset , \U886/U1128/nb , \U886/U1128/na , 
        \U886/U1127/n5 , \U886/U1127/n1 , \U886/U1127/n2 , \U886/U1127/n3 , 
        \U886/U1127/n4 , \U886/U1118_0_/nr , \U886/U1118_0_/nd , 
        \U886/U1118_0_/n2 , \U886/U1118_1_/nr , \U886/U1118_1_/nd , 
        \U886/U1118_1_/n2 , \U886/U1118_2_/nr , \U886/U1118_2_/nd , 
        \U886/U1118_2_/n2 , \U886/U1118_3_/nr , \U886/U1118_3_/nd , 
        \U886/U1118_3_/n2 , \U886/U1117_0_/nr , \U886/U1117_0_/nd , 
        \U886/U1117_0_/n2 , \U886/U1117_1_/nr , \U886/U1117_1_/nd , 
        \U886/U1117_1_/n2 , \U886/U1117_2_/nr , \U886/U1117_2_/nd , 
        \U886/U1117_2_/n2 , \U886/U1117_3_/nr , \U886/U1117_3_/nd , 
        \U886/U1117_3_/n2 , \U884/nack , \U884/acka , \U884/ackb , 
        \U884/reset , \U884/U1128/nb , \U884/U1128/na , \U884/U1127/n5 , 
        \U884/U1127/n1 , \U884/U1127/n2 , \U884/U1127/n3 , \U884/U1127/n4 , 
        \U884/U1118_0_/nr , \U884/U1118_0_/nd , \U884/U1118_0_/n2 , 
        \U884/U1118_1_/nr , \U884/U1118_1_/nd , \U884/U1118_1_/n2 , 
        \U884/U1118_2_/nr , \U884/U1118_2_/nd , \U884/U1118_2_/n2 , 
        \U884/U1118_3_/nr , \U884/U1118_3_/nd , \U884/U1118_3_/n2 , 
        \U884/U1117_0_/nr , \U884/U1117_0_/nd , \U884/U1117_0_/n2 , 
        \U884/U1117_1_/nr , \U884/U1117_1_/nd , \U884/U1117_1_/n2 , 
        \U884/U1117_2_/nr , \U884/U1117_2_/nd , \U884/U1117_2_/n2 , 
        \U884/U1117_3_/nr , \U884/U1117_3_/nd , \U884/U1117_3_/n2 , 
        \U888/naack , \U888/r , \U888/s , \U888/nback , \U888/reset , 
        \U887/naack , \U887/r , \U887/s , \U887/nback , \U887/reset , 
        \U885/naack , \U885/r , \U885/s , \U885/nback , \U885/reset , \U877/x , 
        \U877/y , \U877/reset , \U877/U590/U25/U1/clr , \U877/U590/U25/U1/ob , 
        \U877/U589/U25/U1/clr , \U877/U589/U25/U1/ob , \U877/U588/U25/U1/clr , 
        \U877/U588/U25/U1/ob , \U877/U591/U25/U1/clr , \U877/U591/U25/U1/ob , 
        \U876/x , \U876/y , \U876/reset , \U876/U590/U25/U1/clr , 
        \U876/U590/U25/U1/ob , \U876/U589/U25/U1/clr , \U876/U589/U25/U1/ob , 
        \U876/U588/U25/U1/clr , \U876/U588/U25/U1/ob , \U876/U591/U25/U1/clr , 
        \U876/U591/U25/U1/ob , \U2/x , \U2/y , \U2/reset , 
        \U2/U590/U25/U1/clr , \U2/U590/U25/U1/ob , \U2/U589/U25/U1/clr , 
        \U2/U589/U25/U1/ob , \U2/U588/U25/U1/clr , \U2/U588/U25/U1/ob , 
        \U2/U591/U25/U1/clr , \U2/U591/U25/U1/ob , \U1/x , \U1/y , \U1/reset , 
        \U1/U590/U25/U1/clr , \U1/U590/U25/U1/ob , \U1/U589/U25/U1/clr , 
        \U1/U589/U25/U1/ob , \U1/U588/U25/U1/clr , \U1/U588/U25/U1/ob , 
        \U1/U591/U25/U1/clr , \U1/U591/U25/U1/ob , \U881/nack[1] , 
        \U881/nack[0] , n1;
    buf_2 U897 ( .x(nbReset), .a(nReset) );
    and4_1 \U894/U12  ( .x(eop), .a(ncla), .b(csela), .c(asela), .d(i[4]) );
    inv_1 \U891/U1126/U3  ( .x(\U891/reset ), .a(nbReset) );
    inv_1 \U891/U1139/U3  ( .x(\U891/neopack ), .a(eop) );
    nand3_1 \U891/U1131/U9  ( .x(\U891/iay ), .a(\U891/neopack ), .b(
        \U891/naack[0] ), .c(\U891/naack[1] ) );
    nor3_1 \U891/U1128/U27  ( .x(\U891/U1128/nb ), .a(\U891/reset ), .b(\b[3] 
        ), .c(\b[2] ) );
    nor2_1 \U891/U1128/U26  ( .x(\U891/U1128/na ), .a(\b[1] ), .b(\b[0] ) );
    nand2_2 \U891/U1128/U29  ( .x(\U891/ackb ), .a(\U891/U1128/nb ), .b(
        \U891/U1128/na ) );
    nor2_1 \U891/U1133/U5  ( .x(\U891/naack[0] ), .a(\a[3] ), .b(\a[2] ) );
    nor2_1 \U891/U1108/U5  ( .x(\U891/nack ), .a(\U891/acka ), .b(\U891/ackb )
         );
    nor2_1 \U891/U1134/U5  ( .x(\U891/naack[1] ), .a(\a[1] ), .b(\a[0] ) );
    nor2_2 \U891/U914/U6  ( .x(nia), .a(\U891/iay ), .b(\U891/ackb ) );
    nand2_1 \U891/U1130/U5  ( .x(\U891/acka ), .a(\U891/naack[0] ), .b(
        \U891/naack[1] ) );
    ao222_4 \U891/U1121/U1/U1  ( .x(bsela), .a(\U891/nack ), .b(bsel), .c(
        \U891/nack ), .d(bsela), .e(bsel), .f(bsela) );
    ao222_4 \U891/U1120/U1/U1  ( .x(asela), .a(asel), .b(\U891/nack ), .c(asel
        ), .d(asela), .e(\U891/nack ), .f(asela) );
    nor3_1 \U891/U1118_0_/Unr  ( .x(\U891/U1118_0_/nr ), .a(i[0]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_0_/Und  ( .x(\U891/U1118_0_/nd ), .a(i[0]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_0_/U1  ( .x(\U891/U1118_0_/n2 ), .a(\U891/U1118_0_/n2 ), 
        .b(\U891/U1118_0_/nr ), .c(\U891/U1118_0_/nd ) );
    inv_2 \U891/U1118_0_/U3  ( .x(\a[0] ), .a(\U891/U1118_0_/n2 ) );
    nor3_1 \U891/U1118_1_/Unr  ( .x(\U891/U1118_1_/nr ), .a(i[1]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_1_/Und  ( .x(\U891/U1118_1_/nd ), .a(i[1]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_1_/U1  ( .x(\U891/U1118_1_/n2 ), .a(\U891/U1118_1_/n2 ), 
        .b(\U891/U1118_1_/nr ), .c(\U891/U1118_1_/nd ) );
    inv_2 \U891/U1118_1_/U3  ( .x(\a[1] ), .a(\U891/U1118_1_/n2 ) );
    nor3_1 \U891/U1118_2_/Unr  ( .x(\U891/U1118_2_/nr ), .a(i[2]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_2_/Und  ( .x(\U891/U1118_2_/nd ), .a(i[2]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_2_/U1  ( .x(\U891/U1118_2_/n2 ), .a(\U891/U1118_2_/n2 ), 
        .b(\U891/U1118_2_/nr ), .c(\U891/U1118_2_/nd ) );
    inv_2 \U891/U1118_2_/U3  ( .x(\a[2] ), .a(\U891/U1118_2_/n2 ) );
    nor3_1 \U891/U1118_3_/Unr  ( .x(\U891/U1118_3_/nr ), .a(i[3]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_3_/Und  ( .x(\U891/U1118_3_/nd ), .a(i[3]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_3_/U1  ( .x(\U891/U1118_3_/n2 ), .a(\U891/U1118_3_/n2 ), 
        .b(\U891/U1118_3_/nr ), .c(\U891/U1118_3_/nd ) );
    inv_2 \U891/U1118_3_/U3  ( .x(\a[3] ), .a(\U891/U1118_3_/n2 ) );
    nor3_1 \U891/U1117_0_/Unr  ( .x(\U891/U1117_0_/nr ), .a(i[0]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_0_/Und  ( .x(\U891/U1117_0_/nd ), .a(i[0]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_0_/U1  ( .x(\U891/U1117_0_/n2 ), .a(\U891/U1117_0_/n2 ), 
        .b(\U891/U1117_0_/nr ), .c(\U891/U1117_0_/nd ) );
    inv_2 \U891/U1117_0_/U3  ( .x(\b[0] ), .a(\U891/U1117_0_/n2 ) );
    nor3_1 \U891/U1117_1_/Unr  ( .x(\U891/U1117_1_/nr ), .a(i[1]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_1_/Und  ( .x(\U891/U1117_1_/nd ), .a(i[1]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_1_/U1  ( .x(\U891/U1117_1_/n2 ), .a(\U891/U1117_1_/n2 ), 
        .b(\U891/U1117_1_/nr ), .c(\U891/U1117_1_/nd ) );
    inv_2 \U891/U1117_1_/U3  ( .x(\b[1] ), .a(\U891/U1117_1_/n2 ) );
    nor3_1 \U891/U1117_2_/Unr  ( .x(\U891/U1117_2_/nr ), .a(i[2]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_2_/Und  ( .x(\U891/U1117_2_/nd ), .a(i[2]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_2_/U1  ( .x(\U891/U1117_2_/n2 ), .a(\U891/U1117_2_/n2 ), 
        .b(\U891/U1117_2_/nr ), .c(\U891/U1117_2_/nd ) );
    inv_2 \U891/U1117_2_/U3  ( .x(\b[2] ), .a(\U891/U1117_2_/n2 ) );
    nor3_1 \U891/U1117_3_/Unr  ( .x(\U891/U1117_3_/nr ), .a(i[3]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_3_/Und  ( .x(\U891/U1117_3_/nd ), .a(i[3]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_3_/U1  ( .x(\U891/U1117_3_/n2 ), .a(\U891/U1117_3_/n2 ), 
        .b(\U891/U1117_3_/nr ), .c(\U891/U1117_3_/nd ) );
    inv_2 \U891/U1117_3_/U3  ( .x(\b[3] ), .a(\U891/U1117_3_/n2 ) );
    inv_1 \U886/U1126/U3  ( .x(\U886/reset ), .a(nbReset) );
    nor3_1 \U886/U1128/U27  ( .x(\U886/U1128/nb ), .a(\U886/reset ), .b(\f[3] 
        ), .c(\f[2] ) );
    nor2_1 \U886/U1128/U26  ( .x(\U886/U1128/na ), .a(\f[1] ), .b(\f[0] ) );
    nand2_2 \U886/U1128/U29  ( .x(\U886/ackb ), .a(\U886/U1128/nb ), .b(
        \U886/U1128/na ) );
    nor2_1 \U886/U1108/U5  ( .x(\U886/nack ), .a(\U886/acka ), .b(\U886/ackb )
         );
    nor2_2 \U886/U914/U6  ( .x(nba), .a(\U886/acka ), .b(\U886/ackb ) );
    and4_1 \U886/U1127/U25  ( .x(\U886/U1127/n5 ), .a(\U886/U1127/n1 ), .b(
        \U886/U1127/n2 ), .c(\U886/U1127/n3 ), .d(\U886/U1127/n4 ) );
    inv_1 \U886/U1127/U1  ( .x(\U886/U1127/n1 ), .a(\e[3] ) );
    inv_1 \U886/U1127/U2  ( .x(\U886/U1127/n2 ), .a(\e[2] ) );
    inv_1 \U886/U1127/U3  ( .x(\U886/U1127/n3 ), .a(\e[1] ) );
    inv_1 \U886/U1127/U4  ( .x(\U886/U1127/n4 ), .a(\e[0] ) );
    inv_2 \U886/U1127/U5  ( .x(\U886/acka ), .a(\U886/U1127/n5 ) );
    ao222_2 \U886/U1121/U19/U1/U1  ( .x(fsela), .a(\U886/nack ), .b(fsel), .c(
        \U886/nack ), .d(fsela), .e(fsel), .f(fsela) );
    ao222_2 \U886/U1120/U19/U1/U1  ( .x(esela), .a(esel), .b(\U886/nack ), .c(
        esel), .d(esela), .e(\U886/nack ), .f(esela) );
    nor3_1 \U886/U1118_0_/Unr  ( .x(\U886/U1118_0_/nr ), .a(\b[0] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_0_/Und  ( .x(\U886/U1118_0_/nd ), .a(\b[0] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_0_/U1  ( .x(\U886/U1118_0_/n2 ), .a(\U886/U1118_0_/n2 ), 
        .b(\U886/U1118_0_/nr ), .c(\U886/U1118_0_/nd ) );
    inv_2 \U886/U1118_0_/U3  ( .x(\e[0] ), .a(\U886/U1118_0_/n2 ) );
    nor3_1 \U886/U1118_1_/Unr  ( .x(\U886/U1118_1_/nr ), .a(\b[1] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_1_/Und  ( .x(\U886/U1118_1_/nd ), .a(\b[1] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_1_/U1  ( .x(\U886/U1118_1_/n2 ), .a(\U886/U1118_1_/n2 ), 
        .b(\U886/U1118_1_/nr ), .c(\U886/U1118_1_/nd ) );
    inv_2 \U886/U1118_1_/U3  ( .x(\e[1] ), .a(\U886/U1118_1_/n2 ) );
    nor3_1 \U886/U1118_2_/Unr  ( .x(\U886/U1118_2_/nr ), .a(\b[2] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_2_/Und  ( .x(\U886/U1118_2_/nd ), .a(\b[2] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_2_/U1  ( .x(\U886/U1118_2_/n2 ), .a(\U886/U1118_2_/n2 ), 
        .b(\U886/U1118_2_/nr ), .c(\U886/U1118_2_/nd ) );
    inv_2 \U886/U1118_2_/U3  ( .x(\e[2] ), .a(\U886/U1118_2_/n2 ) );
    nor3_1 \U886/U1118_3_/Unr  ( .x(\U886/U1118_3_/nr ), .a(\b[3] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_3_/Und  ( .x(\U886/U1118_3_/nd ), .a(\b[3] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_3_/U1  ( .x(\U886/U1118_3_/n2 ), .a(\U886/U1118_3_/n2 ), 
        .b(\U886/U1118_3_/nr ), .c(\U886/U1118_3_/nd ) );
    inv_2 \U886/U1118_3_/U3  ( .x(\e[3] ), .a(\U886/U1118_3_/n2 ) );
    nor3_1 \U886/U1117_0_/Unr  ( .x(\U886/U1117_0_/nr ), .a(\b[0] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_0_/Und  ( .x(\U886/U1117_0_/nd ), .a(\b[0] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_0_/U1  ( .x(\U886/U1117_0_/n2 ), .a(\U886/U1117_0_/n2 ), 
        .b(\U886/U1117_0_/nr ), .c(\U886/U1117_0_/nd ) );
    inv_2 \U886/U1117_0_/U3  ( .x(\f[0] ), .a(\U886/U1117_0_/n2 ) );
    nor3_1 \U886/U1117_1_/Unr  ( .x(\U886/U1117_1_/nr ), .a(\b[1] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_1_/Und  ( .x(\U886/U1117_1_/nd ), .a(\b[1] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_1_/U1  ( .x(\U886/U1117_1_/n2 ), .a(\U886/U1117_1_/n2 ), 
        .b(\U886/U1117_1_/nr ), .c(\U886/U1117_1_/nd ) );
    inv_2 \U886/U1117_1_/U3  ( .x(\f[1] ), .a(\U886/U1117_1_/n2 ) );
    nor3_1 \U886/U1117_2_/Unr  ( .x(\U886/U1117_2_/nr ), .a(\b[2] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_2_/Und  ( .x(\U886/U1117_2_/nd ), .a(\b[2] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_2_/U1  ( .x(\U886/U1117_2_/n2 ), .a(\U886/U1117_2_/n2 ), 
        .b(\U886/U1117_2_/nr ), .c(\U886/U1117_2_/nd ) );
    inv_2 \U886/U1117_2_/U3  ( .x(\f[2] ), .a(\U886/U1117_2_/n2 ) );
    nor3_1 \U886/U1117_3_/Unr  ( .x(\U886/U1117_3_/nr ), .a(\b[3] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_3_/Und  ( .x(\U886/U1117_3_/nd ), .a(\b[3] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_3_/U1  ( .x(\U886/U1117_3_/n2 ), .a(\U886/U1117_3_/n2 ), 
        .b(\U886/U1117_3_/nr ), .c(\U886/U1117_3_/nd ) );
    inv_2 \U886/U1117_3_/U3  ( .x(\f[3] ), .a(\U886/U1117_3_/n2 ) );
    inv_1 \U884/U1126/U3  ( .x(\U884/reset ), .a(nbReset) );
    nor3_1 \U884/U1128/U27  ( .x(\U884/U1128/nb ), .a(\U884/reset ), .b(\d[3] 
        ), .c(\d[2] ) );
    nor2_1 \U884/U1128/U26  ( .x(\U884/U1128/na ), .a(\d[1] ), .b(\d[0] ) );
    nand2_2 \U884/U1128/U29  ( .x(\U884/ackb ), .a(\U884/U1128/nb ), .b(
        \U884/U1128/na ) );
    nor2_1 \U884/U1108/U5  ( .x(\U884/nack ), .a(\U884/acka ), .b(\U884/ackb )
         );
    nor2_2 \U884/U914/U6  ( .x(naa), .a(\U884/acka ), .b(\U884/ackb ) );
    and4_1 \U884/U1127/U25  ( .x(\U884/U1127/n5 ), .a(\U884/U1127/n1 ), .b(
        \U884/U1127/n2 ), .c(\U884/U1127/n3 ), .d(\U884/U1127/n4 ) );
    inv_1 \U884/U1127/U1  ( .x(\U884/U1127/n1 ), .a(\c[3] ) );
    inv_1 \U884/U1127/U2  ( .x(\U884/U1127/n2 ), .a(\c[2] ) );
    inv_1 \U884/U1127/U3  ( .x(\U884/U1127/n3 ), .a(\c[1] ) );
    inv_1 \U884/U1127/U4  ( .x(\U884/U1127/n4 ), .a(\c[0] ) );
    inv_2 \U884/U1127/U5  ( .x(\U884/acka ), .a(\U884/U1127/n5 ) );
    ao222_2 \U884/U1121/U19/U1/U1  ( .x(dsela), .a(\U884/nack ), .b(dsel), .c(
        \U884/nack ), .d(dsela), .e(dsel), .f(dsela) );
    ao222_2 \U884/U1120/U19/U1/U1  ( .x(csela), .a(csel), .b(\U884/nack ), .c(
        csel), .d(csela), .e(\U884/nack ), .f(csela) );
    nor3_1 \U884/U1118_0_/Unr  ( .x(\U884/U1118_0_/nr ), .a(\a[0] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_0_/Und  ( .x(\U884/U1118_0_/nd ), .a(\a[0] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_0_/U1  ( .x(\U884/U1118_0_/n2 ), .a(\U884/U1118_0_/n2 ), 
        .b(\U884/U1118_0_/nr ), .c(\U884/U1118_0_/nd ) );
    inv_2 \U884/U1118_0_/U3  ( .x(\c[0] ), .a(\U884/U1118_0_/n2 ) );
    nor3_1 \U884/U1118_1_/Unr  ( .x(\U884/U1118_1_/nr ), .a(\a[1] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_1_/Und  ( .x(\U884/U1118_1_/nd ), .a(\a[1] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_1_/U1  ( .x(\U884/U1118_1_/n2 ), .a(\U884/U1118_1_/n2 ), 
        .b(\U884/U1118_1_/nr ), .c(\U884/U1118_1_/nd ) );
    inv_2 \U884/U1118_1_/U3  ( .x(\c[1] ), .a(\U884/U1118_1_/n2 ) );
    nor3_1 \U884/U1118_2_/Unr  ( .x(\U884/U1118_2_/nr ), .a(\a[2] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_2_/Und  ( .x(\U884/U1118_2_/nd ), .a(\a[2] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_2_/U1  ( .x(\U884/U1118_2_/n2 ), .a(\U884/U1118_2_/n2 ), 
        .b(\U884/U1118_2_/nr ), .c(\U884/U1118_2_/nd ) );
    inv_2 \U884/U1118_2_/U3  ( .x(\c[2] ), .a(\U884/U1118_2_/n2 ) );
    nor3_1 \U884/U1118_3_/Unr  ( .x(\U884/U1118_3_/nr ), .a(\a[3] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_3_/Und  ( .x(\U884/U1118_3_/nd ), .a(\a[3] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_3_/U1  ( .x(\U884/U1118_3_/n2 ), .a(\U884/U1118_3_/n2 ), 
        .b(\U884/U1118_3_/nr ), .c(\U884/U1118_3_/nd ) );
    inv_2 \U884/U1118_3_/U3  ( .x(\c[3] ), .a(\U884/U1118_3_/n2 ) );
    nor3_1 \U884/U1117_0_/Unr  ( .x(\U884/U1117_0_/nr ), .a(\a[0] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_0_/Und  ( .x(\U884/U1117_0_/nd ), .a(\a[0] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_0_/U1  ( .x(\U884/U1117_0_/n2 ), .a(\U884/U1117_0_/n2 ), 
        .b(\U884/U1117_0_/nr ), .c(\U884/U1117_0_/nd ) );
    inv_2 \U884/U1117_0_/U3  ( .x(\d[0] ), .a(\U884/U1117_0_/n2 ) );
    nor3_1 \U884/U1117_1_/Unr  ( .x(\U884/U1117_1_/nr ), .a(\a[1] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_1_/Und  ( .x(\U884/U1117_1_/nd ), .a(\a[1] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_1_/U1  ( .x(\U884/U1117_1_/n2 ), .a(\U884/U1117_1_/n2 ), 
        .b(\U884/U1117_1_/nr ), .c(\U884/U1117_1_/nd ) );
    inv_2 \U884/U1117_1_/U3  ( .x(\d[1] ), .a(\U884/U1117_1_/n2 ) );
    nor3_1 \U884/U1117_2_/Unr  ( .x(\U884/U1117_2_/nr ), .a(\a[2] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_2_/Und  ( .x(\U884/U1117_2_/nd ), .a(\a[2] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_2_/U1  ( .x(\U884/U1117_2_/n2 ), .a(\U884/U1117_2_/n2 ), 
        .b(\U884/U1117_2_/nr ), .c(\U884/U1117_2_/nd ) );
    inv_2 \U884/U1117_2_/U3  ( .x(\d[2] ), .a(\U884/U1117_2_/n2 ) );
    nor3_1 \U884/U1117_3_/Unr  ( .x(\U884/U1117_3_/nr ), .a(\a[3] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_3_/Und  ( .x(\U884/U1117_3_/nd ), .a(\a[3] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_3_/U1  ( .x(\U884/U1117_3_/n2 ), .a(\U884/U1117_3_/n2 ), 
        .b(\U884/U1117_3_/nr ), .c(\U884/U1117_3_/nd ) );
    inv_2 \U884/U1117_3_/U3  ( .x(\d[3] ), .a(\U884/U1117_3_/n2 ) );
    nand2_1 \U888/U1128/U5  ( .x(\U888/s ), .a(\U888/r ), .b(\U888/nback ) );
    nand2_1 \U888/U1103/U5  ( .x(\U888/r ), .a(\U888/naack ), .b(\U888/s ) );
    inv_1 \U888/U1111/U3  ( .x(\U888/reset ), .a(nbReset) );
    inv_1 \U888/U1112/U3  ( .x(\U888/naack ), .a(esela) );
    nor2_1 \U888/U1127/U5  ( .x(\U888/nback ), .a(fsela), .b(\U888/reset ) );
    and2_2 \U888/U1129/U8  ( .x(esel), .a(\U888/nback ), .b(\U888/s ) );
    and2_2 \U888/U1124/U8  ( .x(fsel), .a(\U888/r ), .b(\U888/naack ) );
    nand2_1 \U887/U1128/U5  ( .x(\U887/s ), .a(\U887/r ), .b(\U887/nback ) );
    nand2_1 \U887/U1103/U5  ( .x(\U887/r ), .a(\U887/naack ), .b(\U887/s ) );
    inv_1 \U887/U1111/U3  ( .x(\U887/reset ), .a(nbReset) );
    inv_1 \U887/U1112/U3  ( .x(\U887/naack ), .a(csela) );
    nor2_1 \U887/U1127/U5  ( .x(\U887/nback ), .a(dsela), .b(\U887/reset ) );
    and2_2 \U887/U1129/U8  ( .x(csel), .a(\U887/nback ), .b(\U887/s ) );
    and2_2 \U887/U1124/U8  ( .x(dsel), .a(\U887/r ), .b(\U887/naack ) );
    nand2_1 \U885/U1128/U5  ( .x(\U885/s ), .a(\U885/r ), .b(\U885/nback ) );
    nand2_1 \U885/U1103/U5  ( .x(\U885/r ), .a(\U885/naack ), .b(\U885/s ) );
    inv_1 \U885/U1111/U3  ( .x(\U885/reset ), .a(nbReset) );
    inv_1 \U885/U1112/U3  ( .x(\U885/naack ), .a(asela) );
    nor2_1 \U885/U1127/U5  ( .x(\U885/nback ), .a(bsela), .b(\U885/reset ) );
    and2_2 \U885/U1129/U8  ( .x(asel), .a(\U885/nback ), .b(\U885/s ) );
    and2_2 \U885/U1124/U8  ( .x(bsel), .a(\U885/r ), .b(\U885/naack ) );
    nor3_1 \U877/U594/U7  ( .x(\U877/x ), .a(ol[7]), .b(\U877/reset ), .c(oh
        [7]) );
    nor3_1 \U877/U593/U7  ( .x(\U877/y ), .a(ol[6]), .b(\U877/reset ), .c(oh
        [6]) );
    inv_1 \U877/U604/U3  ( .x(\U877/reset ), .a(nbReset) );
    oa31_1 \U877/U590/U25/U1/Uclr  ( .x(\U877/U590/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[1] ), .d(oh[6]) );
    oaoi211_1 \U877/U590/U25/U1/Uaoi  ( .x(\U877/U590/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[1] ), .c(n1), .d(\U877/U590/U25/U1/clr ) );
    inv_2 \U877/U590/U25/U1/Ui  ( .x(oh[6]), .a(\U877/U590/U25/U1/ob ) );
    oa31_1 \U877/U589/U25/U1/Uclr  ( .x(\U877/U589/U25/U1/clr ), .a(net135), 
        .b(\cl[1] ), .c(\cl[0] ), .d(ol[7]) );
    oaoi211_1 \U877/U589/U25/U1/Uaoi  ( .x(\U877/U589/U25/U1/ob ), .a(\cl[1] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U589/U25/U1/clr ) );
    inv_2 \U877/U589/U25/U1/Ui  ( .x(ol[7]), .a(\U877/U589/U25/U1/ob ) );
    oa31_1 \U877/U588/U25/U1/Uclr  ( .x(\U877/U588/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[2] ), .d(oh[7]) );
    oaoi211_1 \U877/U588/U25/U1/Uaoi  ( .x(\U877/U588/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[2] ), .c(n1), .d(\U877/U588/U25/U1/clr ) );
    inv_2 \U877/U588/U25/U1/Ui  ( .x(oh[7]), .a(\U877/U588/U25/U1/ob ) );
    oa31_1 \U877/U591/U25/U1/Uclr  ( .x(\U877/U591/U25/U1/clr ), .a(net135), 
        .b(\cl[2] ), .c(\cl[0] ), .d(ol[6]) );
    oaoi211_1 \U877/U591/U25/U1/Uaoi  ( .x(\U877/U591/U25/U1/ob ), .a(\cl[2] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U591/U25/U1/clr ) );
    inv_2 \U877/U591/U25/U1/Ui  ( .x(ol[6]), .a(\U877/U591/U25/U1/ob ) );
    ao222_2 \U877/U592/U19/U1/U1  ( .x(ncla), .a(\U877/x ), .b(\U877/y ), .c(
        \U877/x ), .d(ncla), .e(\U877/y ), .f(ncla) );
    nor3_1 \U876/U594/U7  ( .x(\U876/x ), .a(ol[3]), .b(\U876/reset ), .c(oh
        [3]) );
    nor3_1 \U876/U593/U7  ( .x(\U876/y ), .a(ol[2]), .b(\U876/reset ), .c(oh
        [2]) );
    inv_1 \U876/U604/U3  ( .x(\U876/reset ), .a(nbReset) );
    oa31_1 \U876/U590/U25/U1/Uclr  ( .x(\U876/U590/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[1] ), .d(oh[2]) );
    oaoi211_1 \U876/U590/U25/U1/Uaoi  ( .x(\U876/U590/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[1] ), .c(n1), .d(\U876/U590/U25/U1/clr ) );
    inv_2 \U876/U590/U25/U1/Ui  ( .x(oh[2]), .a(\U876/U590/U25/U1/ob ) );
    oa31_1 \U876/U589/U25/U1/Uclr  ( .x(\U876/U589/U25/U1/clr ), .a(net135), 
        .b(\d[1] ), .c(\d[0] ), .d(ol[3]) );
    oaoi211_1 \U876/U589/U25/U1/Uaoi  ( .x(\U876/U589/U25/U1/ob ), .a(\d[1] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U589/U25/U1/clr ) );
    inv_2 \U876/U589/U25/U1/Ui  ( .x(ol[3]), .a(\U876/U589/U25/U1/ob ) );
    oa31_1 \U876/U588/U25/U1/Uclr  ( .x(\U876/U588/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[2] ), .d(oh[3]) );
    oaoi211_1 \U876/U588/U25/U1/Uaoi  ( .x(\U876/U588/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[2] ), .c(n1), .d(\U876/U588/U25/U1/clr ) );
    inv_2 \U876/U588/U25/U1/Ui  ( .x(oh[3]), .a(\U876/U588/U25/U1/ob ) );
    oa31_1 \U876/U591/U25/U1/Uclr  ( .x(\U876/U591/U25/U1/clr ), .a(net135), 
        .b(\d[2] ), .c(\d[0] ), .d(ol[2]) );
    oaoi211_1 \U876/U591/U25/U1/Uaoi  ( .x(\U876/U591/U25/U1/ob ), .a(\d[2] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U591/U25/U1/clr ) );
    inv_2 \U876/U591/U25/U1/Ui  ( .x(ol[2]), .a(\U876/U591/U25/U1/ob ) );
    ao222_2 \U876/U592/U19/U1/U1  ( .x(nda), .a(\U876/x ), .b(\U876/y ), .c(
        \U876/x ), .d(nda), .e(\U876/y ), .f(nda) );
    nor3_1 \U2/U594/U7  ( .x(\U2/x ), .a(ol[1]), .b(\U2/reset ), .c(oh[1]) );
    nor3_1 \U2/U593/U7  ( .x(\U2/y ), .a(ol[0]), .b(\U2/reset ), .c(oh[0]) );
    inv_1 \U2/U604/U3  ( .x(\U2/reset ), .a(nbReset) );
    oa31_1 \U2/U590/U25/U1/Uclr  ( .x(\U2/U590/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[1] ), .d(oh[0]) );
    oaoi211_1 \U2/U590/U25/U1/Uaoi  ( .x(\U2/U590/U25/U1/ob ), .a(\f[3] ), .b(
        \f[1] ), .c(n1), .d(\U2/U590/U25/U1/clr ) );
    inv_2 \U2/U590/U25/U1/Ui  ( .x(oh[0]), .a(\U2/U590/U25/U1/ob ) );
    oa31_1 \U2/U589/U25/U1/Uclr  ( .x(\U2/U589/U25/U1/clr ), .a(net135), .b(
        \f[1] ), .c(\f[0] ), .d(ol[1]) );
    oaoi211_1 \U2/U589/U25/U1/Uaoi  ( .x(\U2/U589/U25/U1/ob ), .a(\f[1] ), .b(
        \f[0] ), .c(n1), .d(\U2/U589/U25/U1/clr ) );
    inv_2 \U2/U589/U25/U1/Ui  ( .x(ol[1]), .a(\U2/U589/U25/U1/ob ) );
    oa31_1 \U2/U588/U25/U1/Uclr  ( .x(\U2/U588/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[2] ), .d(oh[1]) );
    oaoi211_1 \U2/U588/U25/U1/Uaoi  ( .x(\U2/U588/U25/U1/ob ), .a(\f[3] ), .b(
        \f[2] ), .c(n1), .d(\U2/U588/U25/U1/clr ) );
    inv_2 \U2/U588/U25/U1/Ui  ( .x(oh[1]), .a(\U2/U588/U25/U1/ob ) );
    oa31_1 \U2/U591/U25/U1/Uclr  ( .x(\U2/U591/U25/U1/clr ), .a(net135), .b(
        \f[2] ), .c(\f[0] ), .d(ol[0]) );
    oaoi211_1 \U2/U591/U25/U1/Uaoi  ( .x(\U2/U591/U25/U1/ob ), .a(\f[2] ), .b(
        \f[0] ), .c(n1), .d(\U2/U591/U25/U1/clr ) );
    inv_2 \U2/U591/U25/U1/Ui  ( .x(ol[0]), .a(\U2/U591/U25/U1/ob ) );
    ao222_2 \U2/U592/U19/U1/U1  ( .x(nfa), .a(\U2/x ), .b(\U2/y ), .c(\U2/x ), 
        .d(nfa), .e(\U2/y ), .f(nfa) );
    nor3_1 \U1/U594/U7  ( .x(\U1/x ), .a(ol[5]), .b(\U1/reset ), .c(oh[5]) );
    nor3_1 \U1/U593/U7  ( .x(\U1/y ), .a(ol[4]), .b(\U1/reset ), .c(oh[4]) );
    inv_1 \U1/U604/U3  ( .x(\U1/reset ), .a(nbReset) );
    oa31_1 \U1/U590/U25/U1/Uclr  ( .x(\U1/U590/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[1] ), .d(oh[4]) );
    oaoi211_1 \U1/U590/U25/U1/Uaoi  ( .x(\U1/U590/U25/U1/ob ), .a(\e[3] ), .b(
        \e[1] ), .c(n1), .d(\U1/U590/U25/U1/clr ) );
    inv_2 \U1/U590/U25/U1/Ui  ( .x(oh[4]), .a(\U1/U590/U25/U1/ob ) );
    oa31_1 \U1/U589/U25/U1/Uclr  ( .x(\U1/U589/U25/U1/clr ), .a(net135), .b(
        \e[1] ), .c(\e[0] ), .d(ol[5]) );
    oaoi211_1 \U1/U589/U25/U1/Uaoi  ( .x(\U1/U589/U25/U1/ob ), .a(\e[1] ), .b(
        \e[0] ), .c(n1), .d(\U1/U589/U25/U1/clr ) );
    inv_2 \U1/U589/U25/U1/Ui  ( .x(ol[5]), .a(\U1/U589/U25/U1/ob ) );
    oa31_1 \U1/U588/U25/U1/Uclr  ( .x(\U1/U588/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[2] ), .d(oh[5]) );
    oaoi211_1 \U1/U588/U25/U1/Uaoi  ( .x(\U1/U588/U25/U1/ob ), .a(\e[3] ), .b(
        \e[2] ), .c(n1), .d(\U1/U588/U25/U1/clr ) );
    inv_2 \U1/U588/U25/U1/Ui  ( .x(oh[5]), .a(\U1/U588/U25/U1/ob ) );
    oa31_1 \U1/U591/U25/U1/Uclr  ( .x(\U1/U591/U25/U1/clr ), .a(net135), .b(
        \e[2] ), .c(\e[0] ), .d(ol[4]) );
    oaoi211_1 \U1/U591/U25/U1/Uaoi  ( .x(\U1/U591/U25/U1/ob ), .a(\e[2] ), .b(
        \e[0] ), .c(n1), .d(\U1/U591/U25/U1/clr ) );
    inv_2 \U1/U591/U25/U1/Ui  ( .x(ol[4]), .a(\U1/U591/U25/U1/ob ) );
    ao222_2 \U1/U592/U19/U1/U1  ( .x(nea), .a(\U1/x ), .b(\U1/y ), .c(\U1/x ), 
        .d(nea), .e(\U1/y ), .f(nea) );
    and3_4 \U881/U20/U9  ( .x(nca), .a(\U881/nack[1] ), .b(\U881/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U881/U18/U5  ( .x(\U881/nack[0] ), .a(\cl[3] ), .b(\cl[0] ) );
    nor2_1 \U881/U19/U5  ( .x(\U881/nack[1] ), .a(\cl[1] ), .b(\cl[2] ) );
    ao222_2 \U881/U15_0_/U19/U1/U1  ( .x(\cl[0] ), .a(\c[0] ), .b(ncla), .c(
        \c[0] ), .d(\cl[0] ), .e(ncla), .f(\cl[0] ) );
    ao222_2 \U881/U15_1_/U19/U1/U1  ( .x(\cl[1] ), .a(\c[1] ), .b(ncla), .c(
        \c[1] ), .d(\cl[1] ), .e(ncla), .f(\cl[1] ) );
    ao222_2 \U881/U15_2_/U19/U1/U1  ( .x(\cl[2] ), .a(\c[2] ), .b(ncla), .c(
        \c[2] ), .d(\cl[2] ), .e(ncla), .f(\cl[2] ) );
    ao222_2 \U881/U15_3_/U19/U1/U1  ( .x(\cl[3] ), .a(\c[3] ), .b(ncla), .c(
        \c[3] ), .d(\cl[3] ), .e(ncla), .f(\cl[3] ) );
    and2_5 U1 ( .x(n1), .a(nbReset), .b(noa) );
    and2_3 U2 ( .x(net135), .a(nbReset), .b(noa) );
endmodule


module chain_dr2fr_byte_0 ( eop_ack, ia, o, eop, ih, il, nReset, noa );
output [4:0] o;
input  [7:0] ih;
input  [7:0] il;
input  eop, nReset, noa;
output eop_ack, ia;
    wire eop_pass, nhighack, nlowack, \twobitack[2] , \twobitack[3] , 
        \twobitack[0] , \twobitack[1] , xsel, ysel, nxa, nyla, nbReset, nya, 
        \y[3] , \y[2] , \y[1] , \y[0] , \yl[3] , \yl[2] , \yl[1] , \yl[0] , 
        \cdh[0] , \cdh[1] , \cdl[0] , \cdl[1] , net193, \cdh[2] , \cdh[3] , 
        \cdl[2] , \cdl[3] , net195, bsel, dsel, nba, bg, nda, dg, asel, csel, 
        naa, ag, nca, cg, \d[3] , \d[2] , \d[1] , \d[0] , \b[3] , \b[2] , 
        \b[1] , \b[0] , \x[3] , \x[2] , \x[1] , \x[0] , \c[3] , \c[2] , \c[1] , 
        \c[0] , \a[3] , \a[2] , \a[1] , \a[0] , net194, net199, \U1018/Z , 
        \U1270/net190 , \U1270/net191 , \U1270/net192 , \U1270/net189 , 
        \U1270/U1141/Z , \U1268/net190 , \U1268/net191 , \U1268/net192 , 
        \U1268/net189 , \U1268/U1141/Z , \U1224/nack[0] , \U1224/nack[1] , 
        \U1224/net4 , \U1224/U1125/U28/U1/clr , \U1224/U1125/U28/U1/set , 
        \U1224/U1122/U28/U1/clr , \U1224/U1122/U28/U1/set , 
        \U1224/U916_0_/U25/U1/clr , \U1224/U916_0_/U25/U1/ob , 
        \U1224/U916_1_/U25/U1/clr , \U1224/U916_1_/U25/U1/ob , 
        \U1224/U916_2_/U25/U1/clr , \U1224/U916_2_/U25/U1/ob , 
        \U1224/U916_3_/U25/U1/clr , \U1224/U916_3_/U25/U1/ob , \U1209/nack[0] , 
        \U1209/nack[1] , \U1209/net4 , \U1209/U1125/U28/U1/clr , 
        \U1209/U1125/U28/U1/set , \U1209/U1122/U28/U1/clr , 
        \U1209/U1122/U28/U1/set , \U1209/U916_0_/U25/U1/clr , 
        \U1209/U916_0_/U25/U1/ob , \U1209/U916_1_/U25/U1/clr , 
        \U1209/U916_1_/U25/U1/ob , \U1209/U916_2_/U25/U1/clr , 
        \U1209/U916_2_/U25/U1/ob , \U1209/U916_3_/U25/U1/clr , 
        \U1209/U916_3_/U25/U1/ob , \U1213/nack[0] , \U1213/nack[1] , 
        \U1213/net4 , \U1213/U1125/U28/U1/clr , \U1213/U1125/U28/U1/set , 
        \U1213/U1122/U28/U1/clr , \U1213/U1122/U28/U1/set , 
        \U1213/U916_0_/U25/U1/clr , \U1213/U916_0_/U25/U1/ob , 
        \U1213/U916_1_/U25/U1/clr , \U1213/U916_1_/U25/U1/ob , 
        \U1213/U916_2_/U25/U1/clr , \U1213/U916_2_/U25/U1/ob , 
        \U1213/U916_3_/U25/U1/clr , \U1213/U916_3_/U25/U1/ob , \U1296/ng , 
        \U1296/U1384/Z , \U1296/U1386/U25/U1/clr , \U1296/U1386/U25/U1/ob , 
        \U1298/ng , \U1298/U1384/Z , \U1298/U1386/U25/U1/clr , 
        \U1298/U1386/U25/U1/ob , \U1306/ng , \U1306/U1384/Z , 
        \U1306/U1386/U25/U1/clr , \U1306/U1386/U25/U1/ob , \U1295/ng , 
        \U1295/U1384/Z , \U1295/U1386/U25/U1/clr , \U1295/U1386/U25/U1/ob , 
        \U1297/s , \U1297/nback , \U1297/r , \U1297/naack , \U1297/reset , 
        \U1297/U1128/U28/U1/clr , \U1297/U1128/U28/U1/set , 
        \U1297/U1127/U28/U1/clr , \U1297/U1127/U28/U1/set , \U1300/s , 
        \U1300/nback , \U1300/r , \U1300/naack , \U1300/reset , 
        \U1300/U1128/U28/U1/clr , \U1300/U1128/U28/U1/set , 
        \U1300/U1127/U28/U1/clr , \U1300/U1127/U28/U1/set , \U1289/bnreset , 
        \U1289/U1150/U28/U1/clr , \U1289/U1150/U28/U1/set , 
        \U1289/U1152/U28/U1/clr , \U1289/U1152/U28/U1/set , 
        \U1289/U1149/U28/U1/clr , \U1289/U1149/U28/U1/set , 
        \U1289/U1151/U28/U1/clr , \U1289/U1151/U28/U1/set , 
        \U1289/U1148/net190 , \U1289/U1148/net191 , \U1289/U1148/net192 , 
        \U1289/U1148/net189 , \U1289/U1148/U1141/Z , \U1271/bnreset , 
        \U1271/U1150/U28/U1/clr , \U1271/U1150/U28/U1/set , 
        \U1271/U1152/U28/U1/clr , \U1271/U1152/U28/U1/set , 
        \U1271/U1149/U28/U1/clr , \U1271/U1149/U28/U1/set , 
        \U1271/U1151/U28/U1/clr , \U1271/U1151/U28/U1/set , 
        \U1271/U1148/net190 , \U1271/U1148/net191 , \U1271/U1148/net192 , 
        \U1271/U1148/net189 , \U1271/U1148/U1141/Z , \U1225/naack , \U1225/r , 
        \U1225/s , \U1225/nback , \U1225/reset , \U1308/nack[1] , 
        \U1308/nack[0] ;
    assign o[4] = eop_ack;
    buf_2 U1231 ( .x(nbReset), .a(nReset) );
    and3_1 \U1194/U9  ( .x(eop_pass), .a(nxa), .b(naa), .c(eop) );
    ao222_1 \U1301/U18/U1/U1  ( .x(nlowack), .a(\twobitack[0] ), .b(
        \twobitack[1] ), .c(\twobitack[0] ), .d(nlowack), .e(\twobitack[1] ), 
        .f(nlowack) );
    ao222_1 \U1302/U18/U1/U1  ( .x(nhighack), .a(\twobitack[2] ), .b(
        \twobitack[3] ), .c(\twobitack[2] ), .d(nhighack), .e(\twobitack[3] ), 
        .f(nhighack) );
    aoi222_1 \U1018/U30/U1  ( .x(ia), .a(nhighack), .b(nlowack), .c(nhighack), 
        .d(\U1018/Z ), .e(nlowack), .f(\U1018/Z ) );
    inv_1 \U1018/U30/Uinv  ( .x(\U1018/Z ), .a(ia) );
    ao222_2 \U1038/U19/U1/U1  ( .x(eop_ack), .a(eop_pass), .b(noa), .c(
        eop_pass), .d(eop_ack), .e(noa), .f(eop_ack) );
    inv_1 \U1270/U1147/U3  ( .x(\U1270/net189 ), .a(nbReset) );
    nor2_1 \U1270/U582/U5  ( .x(\U1270/net192 ), .a(il[4]), .b(ih[4]) );
    nor2_1 \U1270/U580/U5  ( .x(\U1270/net191 ), .a(il[5]), .b(ih[5]) );
    nor2_2 \U1270/U1146/U6  ( .x(net199), .a(\U1270/net190 ), .b(
        \U1270/net189 ) );
    aoi222_1 \U1270/U1141/U30/U1  ( .x(\U1270/net190 ), .a(\U1270/net191 ), 
        .b(\U1270/net192 ), .c(\U1270/net191 ), .d(\U1270/U1141/Z ), .e(
        \U1270/net192 ), .f(\U1270/U1141/Z ) );
    inv_1 \U1270/U1141/U30/Uinv  ( .x(\U1270/U1141/Z ), .a(\U1270/net190 ) );
    inv_1 \U1268/U1147/U3  ( .x(\U1268/net189 ), .a(nbReset) );
    nor2_1 \U1268/U582/U5  ( .x(\U1268/net192 ), .a(il[6]), .b(ih[6]) );
    nor2_1 \U1268/U580/U5  ( .x(\U1268/net191 ), .a(il[7]), .b(ih[7]) );
    nor2_2 \U1268/U1146/U6  ( .x(net194), .a(\U1268/net190 ), .b(
        \U1268/net189 ) );
    aoi222_1 \U1268/U1141/U30/U1  ( .x(\U1268/net190 ), .a(\U1268/net191 ), 
        .b(\U1268/net192 ), .c(\U1268/net191 ), .d(\U1268/U1141/Z ), .e(
        \U1268/net192 ), .f(\U1268/U1141/Z ) );
    inv_1 \U1268/U1141/U30/Uinv  ( .x(\U1268/U1141/Z ), .a(\U1268/net190 ) );
    nor2_1 \U1224/U1128/U5  ( .x(\U1224/nack[0] ), .a(\x[3] ), .b(\x[2] ) );
    nor3_1 \U1224/U1127/U7  ( .x(\U1224/nack[1] ), .a(\x[1] ), .b(\U1224/net4 
        ), .c(\x[0] ) );
    inv_1 \U1224/U907/U3  ( .x(\U1224/net4 ), .a(nbReset) );
    aoai211_1 \U1224/U1125/U28/U1/U1  ( .x(\U1224/U1125/U28/U1/clr ), .a(
        \U1224/nack[1] ), .b(\U1224/nack[0] ), .c(asel), .d(naa) );
    nand3_1 \U1224/U1125/U28/U1/U2  ( .x(\U1224/U1125/U28/U1/set ), .a(asel), 
        .b(\U1224/nack[1] ), .c(\U1224/nack[0] ) );
    nand2_2 \U1224/U1125/U28/U1/U3  ( .x(naa), .a(\U1224/U1125/U28/U1/clr ), 
        .b(\U1224/U1125/U28/U1/set ) );
    aoai211_1 \U1224/U1122/U28/U1/U1  ( .x(\U1224/U1122/U28/U1/clr ), .a(
        \U1224/nack[0] ), .b(\U1224/nack[1] ), .c(csel), .d(nca) );
    nand3_1 \U1224/U1122/U28/U1/U2  ( .x(\U1224/U1122/U28/U1/set ), .a(csel), 
        .b(\U1224/nack[0] ), .c(\U1224/nack[1] ) );
    nand2_2 \U1224/U1122/U28/U1/U3  ( .x(nca), .a(\U1224/U1122/U28/U1/clr ), 
        .b(\U1224/U1122/U28/U1/set ) );
    oa31_1 \U1224/U916_0_/U25/U1/Uclr  ( .x(\U1224/U916_0_/U25/U1/clr ), .a(
        nxa), .b(\a[0] ), .c(\c[0] ), .d(\x[0] ) );
    oaoi211_1 \U1224/U916_0_/U25/U1/Uaoi  ( .x(\U1224/U916_0_/U25/U1/ob ), .a(
        \a[0] ), .b(\c[0] ), .c(nxa), .d(\U1224/U916_0_/U25/U1/clr ) );
    inv_2 \U1224/U916_0_/U25/U1/Ui  ( .x(\x[0] ), .a(\U1224/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_1_/U25/U1/Uclr  ( .x(\U1224/U916_1_/U25/U1/clr ), .a(
        nxa), .b(\a[1] ), .c(\c[1] ), .d(\x[1] ) );
    oaoi211_1 \U1224/U916_1_/U25/U1/Uaoi  ( .x(\U1224/U916_1_/U25/U1/ob ), .a(
        \a[1] ), .b(\c[1] ), .c(nxa), .d(\U1224/U916_1_/U25/U1/clr ) );
    inv_2 \U1224/U916_1_/U25/U1/Ui  ( .x(\x[1] ), .a(\U1224/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_2_/U25/U1/Uclr  ( .x(\U1224/U916_2_/U25/U1/clr ), .a(
        nxa), .b(\a[2] ), .c(\c[2] ), .d(\x[2] ) );
    oaoi211_1 \U1224/U916_2_/U25/U1/Uaoi  ( .x(\U1224/U916_2_/U25/U1/ob ), .a(
        \a[2] ), .b(\c[2] ), .c(nxa), .d(\U1224/U916_2_/U25/U1/clr ) );
    inv_2 \U1224/U916_2_/U25/U1/Ui  ( .x(\x[2] ), .a(\U1224/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_3_/U25/U1/Uclr  ( .x(\U1224/U916_3_/U25/U1/clr ), .a(
        nxa), .b(\a[3] ), .c(\c[3] ), .d(\x[3] ) );
    oaoi211_1 \U1224/U916_3_/U25/U1/Uaoi  ( .x(\U1224/U916_3_/U25/U1/ob ), .a(
        \a[3] ), .b(\c[3] ), .c(nxa), .d(\U1224/U916_3_/U25/U1/clr ) );
    inv_2 \U1224/U916_3_/U25/U1/Ui  ( .x(\x[3] ), .a(\U1224/U916_3_/U25/U1/ob 
        ) );
    nor2_1 \U1209/U1128/U5  ( .x(\U1209/nack[0] ), .a(o[3]), .b(o[2]) );
    nor3_1 \U1209/U1127/U7  ( .x(\U1209/nack[1] ), .a(o[1]), .b(\U1209/net4 ), 
        .c(o[0]) );
    inv_1 \U1209/U907/U3  ( .x(\U1209/net4 ), .a(nbReset) );
    aoai211_1 \U1209/U1125/U28/U1/U1  ( .x(\U1209/U1125/U28/U1/clr ), .a(
        \U1209/nack[1] ), .b(\U1209/nack[0] ), .c(xsel), .d(nxa) );
    nand3_1 \U1209/U1125/U28/U1/U2  ( .x(\U1209/U1125/U28/U1/set ), .a(xsel), 
        .b(\U1209/nack[1] ), .c(\U1209/nack[0] ) );
    nand2_2 \U1209/U1125/U28/U1/U3  ( .x(nxa), .a(\U1209/U1125/U28/U1/clr ), 
        .b(\U1209/U1125/U28/U1/set ) );
    aoai211_1 \U1209/U1122/U28/U1/U1  ( .x(\U1209/U1122/U28/U1/clr ), .a(
        \U1209/nack[0] ), .b(\U1209/nack[1] ), .c(ysel), .d(nyla) );
    nand3_1 \U1209/U1122/U28/U1/U2  ( .x(\U1209/U1122/U28/U1/set ), .a(ysel), 
        .b(\U1209/nack[0] ), .c(\U1209/nack[1] ) );
    nand2_2 \U1209/U1122/U28/U1/U3  ( .x(nyla), .a(\U1209/U1122/U28/U1/clr ), 
        .b(\U1209/U1122/U28/U1/set ) );
    oa31_1 \U1209/U916_0_/U25/U1/Uclr  ( .x(\U1209/U916_0_/U25/U1/clr ), .a(
        noa), .b(\x[0] ), .c(\yl[0] ), .d(o[0]) );
    oaoi211_1 \U1209/U916_0_/U25/U1/Uaoi  ( .x(\U1209/U916_0_/U25/U1/ob ), .a(
        \x[0] ), .b(\yl[0] ), .c(noa), .d(\U1209/U916_0_/U25/U1/clr ) );
    inv_2 \U1209/U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U1209/U916_0_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_1_/U25/U1/Uclr  ( .x(\U1209/U916_1_/U25/U1/clr ), .a(
        noa), .b(\x[1] ), .c(\yl[1] ), .d(o[1]) );
    oaoi211_1 \U1209/U916_1_/U25/U1/Uaoi  ( .x(\U1209/U916_1_/U25/U1/ob ), .a(
        \x[1] ), .b(\yl[1] ), .c(noa), .d(\U1209/U916_1_/U25/U1/clr ) );
    inv_2 \U1209/U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U1209/U916_1_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_2_/U25/U1/Uclr  ( .x(\U1209/U916_2_/U25/U1/clr ), .a(
        noa), .b(\x[2] ), .c(\yl[2] ), .d(o[2]) );
    oaoi211_1 \U1209/U916_2_/U25/U1/Uaoi  ( .x(\U1209/U916_2_/U25/U1/ob ), .a(
        \x[2] ), .b(\yl[2] ), .c(noa), .d(\U1209/U916_2_/U25/U1/clr ) );
    inv_2 \U1209/U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U1209/U916_2_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_3_/U25/U1/Uclr  ( .x(\U1209/U916_3_/U25/U1/clr ), .a(
        noa), .b(\x[3] ), .c(\yl[3] ), .d(o[3]) );
    oaoi211_1 \U1209/U916_3_/U25/U1/Uaoi  ( .x(\U1209/U916_3_/U25/U1/ob ), .a(
        \x[3] ), .b(\yl[3] ), .c(noa), .d(\U1209/U916_3_/U25/U1/clr ) );
    inv_2 \U1209/U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U1209/U916_3_/U25/U1/ob )
         );
    nor2_1 \U1213/U1128/U5  ( .x(\U1213/nack[0] ), .a(\y[3] ), .b(\y[2] ) );
    nor3_1 \U1213/U1127/U7  ( .x(\U1213/nack[1] ), .a(\y[1] ), .b(\U1213/net4 
        ), .c(\y[0] ) );
    inv_1 \U1213/U907/U3  ( .x(\U1213/net4 ), .a(nbReset) );
    aoai211_1 \U1213/U1125/U28/U1/U1  ( .x(\U1213/U1125/U28/U1/clr ), .a(
        \U1213/nack[1] ), .b(\U1213/nack[0] ), .c(bsel), .d(nba) );
    nand3_1 \U1213/U1125/U28/U1/U2  ( .x(\U1213/U1125/U28/U1/set ), .a(bsel), 
        .b(\U1213/nack[1] ), .c(\U1213/nack[0] ) );
    nand2_2 \U1213/U1125/U28/U1/U3  ( .x(nba), .a(\U1213/U1125/U28/U1/clr ), 
        .b(\U1213/U1125/U28/U1/set ) );
    aoai211_1 \U1213/U1122/U28/U1/U1  ( .x(\U1213/U1122/U28/U1/clr ), .a(
        \U1213/nack[0] ), .b(\U1213/nack[1] ), .c(dsel), .d(nda) );
    nand3_1 \U1213/U1122/U28/U1/U2  ( .x(\U1213/U1122/U28/U1/set ), .a(dsel), 
        .b(\U1213/nack[0] ), .c(\U1213/nack[1] ) );
    nand2_2 \U1213/U1122/U28/U1/U3  ( .x(nda), .a(\U1213/U1122/U28/U1/clr ), 
        .b(\U1213/U1122/U28/U1/set ) );
    oa31_1 \U1213/U916_0_/U25/U1/Uclr  ( .x(\U1213/U916_0_/U25/U1/clr ), .a(
        nya), .b(\b[0] ), .c(\d[0] ), .d(\y[0] ) );
    oaoi211_1 \U1213/U916_0_/U25/U1/Uaoi  ( .x(\U1213/U916_0_/U25/U1/ob ), .a(
        \b[0] ), .b(\d[0] ), .c(nya), .d(\U1213/U916_0_/U25/U1/clr ) );
    inv_2 \U1213/U916_0_/U25/U1/Ui  ( .x(\y[0] ), .a(\U1213/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_1_/U25/U1/Uclr  ( .x(\U1213/U916_1_/U25/U1/clr ), .a(
        nya), .b(\b[1] ), .c(\d[1] ), .d(\y[1] ) );
    oaoi211_1 \U1213/U916_1_/U25/U1/Uaoi  ( .x(\U1213/U916_1_/U25/U1/ob ), .a(
        \b[1] ), .b(\d[1] ), .c(nya), .d(\U1213/U916_1_/U25/U1/clr ) );
    inv_2 \U1213/U916_1_/U25/U1/Ui  ( .x(\y[1] ), .a(\U1213/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_2_/U25/U1/Uclr  ( .x(\U1213/U916_2_/U25/U1/clr ), .a(
        nya), .b(\b[2] ), .c(\d[2] ), .d(\y[2] ) );
    oaoi211_1 \U1213/U916_2_/U25/U1/Uaoi  ( .x(\U1213/U916_2_/U25/U1/ob ), .a(
        \b[2] ), .b(\d[2] ), .c(nya), .d(\U1213/U916_2_/U25/U1/clr ) );
    inv_2 \U1213/U916_2_/U25/U1/Ui  ( .x(\y[2] ), .a(\U1213/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_3_/U25/U1/Uclr  ( .x(\U1213/U916_3_/U25/U1/clr ), .a(
        nya), .b(\b[3] ), .c(\d[3] ), .d(\y[3] ) );
    oaoi211_1 \U1213/U916_3_/U25/U1/Uaoi  ( .x(\U1213/U916_3_/U25/U1/ob ), .a(
        \b[3] ), .b(\d[3] ), .c(nya), .d(\U1213/U916_3_/U25/U1/clr ) );
    inv_2 \U1213/U916_3_/U25/U1/Ui  ( .x(\y[3] ), .a(\U1213/U916_3_/U25/U1/ob 
        ) );
    and3_2 \U1210/U1138/U9  ( .x(\d[3] ), .a(\cdh[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1137/U9  ( .x(\d[2] ), .a(\cdl[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1139/U9  ( .x(\d[1] ), .a(\cdh[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1210/U1136/U9  ( .x(\d[0] ), .a(\cdl[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1162/U1138/U9  ( .x(\a[3] ), .a(ih[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1137/U9  ( .x(\a[2] ), .a(il[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1139/U9  ( .x(\a[1] ), .a(ih[6]), .b(naa), .c(il[7]) );
    and3_2 \U1162/U1136/U9  ( .x(\a[0] ), .a(il[6]), .b(naa), .c(il[7]) );
    and3_2 \U1211/U1138/U9  ( .x(\b[3] ), .a(ih[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1137/U9  ( .x(\b[2] ), .a(il[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1139/U9  ( .x(\b[1] ), .a(ih[4]), .b(nba), .c(il[5]) );
    and3_2 \U1211/U1136/U9  ( .x(\b[0] ), .a(il[4]), .b(nba), .c(il[5]) );
    and3_2 \U1163/U1138/U9  ( .x(\c[3] ), .a(\cdh[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1137/U9  ( .x(\c[2] ), .a(\cdl[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1139/U9  ( .x(\c[1] ), .a(\cdh[2] ), .b(nca), .c(\cdl[3] )
         );
    and3_2 \U1163/U1136/U9  ( .x(\c[0] ), .a(\cdl[2] ), .b(nca), .c(\cdl[3] )
         );
    and2_1 \U1296/U1385/U8  ( .x(cg), .a(nbReset), .b(\U1296/ng ) );
    aoi222_1 \U1296/U1384/U30/U1  ( .x(\U1296/ng ), .a(nca), .b(net195), .c(
        nca), .d(\U1296/U1384/Z ), .e(net195), .f(\U1296/U1384/Z ) );
    inv_1 \U1296/U1384/U30/Uinv  ( .x(\U1296/U1384/Z ), .a(\U1296/ng ) );
    oa31_1 \U1296/U1386/U25/U1/Uclr  ( .x(\U1296/U1386/U25/U1/clr ), .a(
        \twobitack[2] ), .b(cg), .c(nca), .d(net195) );
    oaoi211_1 \U1296/U1386/U25/U1/Uaoi  ( .x(\U1296/U1386/U25/U1/ob ), .a(cg), 
        .b(nca), .c(\twobitack[2] ), .d(\U1296/U1386/U25/U1/clr ) );
    inv_2 \U1296/U1386/U25/U1/Ui  ( .x(net195), .a(\U1296/U1386/U25/U1/ob ) );
    and2_1 \U1298/U1385/U8  ( .x(dg), .a(nbReset), .b(\U1298/ng ) );
    aoi222_1 \U1298/U1384/U30/U1  ( .x(\U1298/ng ), .a(nda), .b(net193), .c(
        nda), .d(\U1298/U1384/Z ), .e(net193), .f(\U1298/U1384/Z ) );
    inv_1 \U1298/U1384/U30/Uinv  ( .x(\U1298/U1384/Z ), .a(\U1298/ng ) );
    oa31_1 \U1298/U1386/U25/U1/Uclr  ( .x(\U1298/U1386/U25/U1/clr ), .a(
        \twobitack[0] ), .b(dg), .c(nda), .d(net193) );
    oaoi211_1 \U1298/U1386/U25/U1/Uaoi  ( .x(\U1298/U1386/U25/U1/ob ), .a(dg), 
        .b(nda), .c(\twobitack[0] ), .d(\U1298/U1386/U25/U1/clr ) );
    inv_2 \U1298/U1386/U25/U1/Ui  ( .x(net193), .a(\U1298/U1386/U25/U1/ob ) );
    and2_1 \U1306/U1385/U8  ( .x(bg), .a(nbReset), .b(\U1306/ng ) );
    aoi222_1 \U1306/U1384/U30/U1  ( .x(\U1306/ng ), .a(nba), .b(\twobitack[1] 
        ), .c(nba), .d(\U1306/U1384/Z ), .e(\twobitack[1] ), .f(
        \U1306/U1384/Z ) );
    inv_1 \U1306/U1384/U30/Uinv  ( .x(\U1306/U1384/Z ), .a(\U1306/ng ) );
    oa31_1 \U1306/U1386/U25/U1/Uclr  ( .x(\U1306/U1386/U25/U1/clr ), .a(net199
        ), .b(bg), .c(nba), .d(\twobitack[1] ) );
    oaoi211_1 \U1306/U1386/U25/U1/Uaoi  ( .x(\U1306/U1386/U25/U1/ob ), .a(bg), 
        .b(nba), .c(net199), .d(\U1306/U1386/U25/U1/clr ) );
    inv_2 \U1306/U1386/U25/U1/Ui  ( .x(\twobitack[1] ), .a(
        \U1306/U1386/U25/U1/ob ) );
    and2_1 \U1295/U1385/U8  ( .x(ag), .a(nbReset), .b(\U1295/ng ) );
    aoi222_1 \U1295/U1384/U30/U1  ( .x(\U1295/ng ), .a(naa), .b(\twobitack[3] 
        ), .c(naa), .d(\U1295/U1384/Z ), .e(\twobitack[3] ), .f(
        \U1295/U1384/Z ) );
    inv_1 \U1295/U1384/U30/Uinv  ( .x(\U1295/U1384/Z ), .a(\U1295/ng ) );
    oa31_1 \U1295/U1386/U25/U1/Uclr  ( .x(\U1295/U1386/U25/U1/clr ), .a(net194
        ), .b(ag), .c(naa), .d(\twobitack[3] ) );
    oaoi211_1 \U1295/U1386/U25/U1/Uaoi  ( .x(\U1295/U1386/U25/U1/ob ), .a(ag), 
        .b(naa), .c(net194), .d(\U1295/U1386/U25/U1/clr ) );
    inv_2 \U1295/U1386/U25/U1/Ui  ( .x(\twobitack[3] ), .a(
        \U1295/U1386/U25/U1/ob ) );
    nand2_1 \U1297/U1131/U5  ( .x(\U1297/s ), .a(\U1297/r ), .b(\U1297/nback )
         );
    nand2_1 \U1297/U1103/U5  ( .x(\U1297/r ), .a(\U1297/naack ), .b(\U1297/s )
         );
    inv_1 \U1297/U1111/U3  ( .x(\U1297/reset ), .a(nbReset) );
    inv_1 \U1297/U1112/U3  ( .x(\U1297/naack ), .a(naa) );
    nor2_1 \U1297/U1130/U5  ( .x(\U1297/nback ), .a(nca), .b(\U1297/reset ) );
    aoai211_1 \U1297/U1128/U28/U1/U1  ( .x(\U1297/U1128/U28/U1/clr ), .a(
        \U1297/r ), .b(\U1297/naack ), .c(cg), .d(csel) );
    nand3_1 \U1297/U1128/U28/U1/U2  ( .x(\U1297/U1128/U28/U1/set ), .a(cg), 
        .b(\U1297/r ), .c(\U1297/naack ) );
    nand2_2 \U1297/U1128/U28/U1/U3  ( .x(csel), .a(\U1297/U1128/U28/U1/clr ), 
        .b(\U1297/U1128/U28/U1/set ) );
    aoai211_1 \U1297/U1127/U28/U1/U1  ( .x(\U1297/U1127/U28/U1/clr ), .a(
        \U1297/s ), .b(\U1297/nback ), .c(ag), .d(asel) );
    nand3_1 \U1297/U1127/U28/U1/U2  ( .x(\U1297/U1127/U28/U1/set ), .a(ag), 
        .b(\U1297/s ), .c(\U1297/nback ) );
    nand2_2 \U1297/U1127/U28/U1/U3  ( .x(asel), .a(\U1297/U1127/U28/U1/clr ), 
        .b(\U1297/U1127/U28/U1/set ) );
    nand2_1 \U1300/U1131/U5  ( .x(\U1300/s ), .a(\U1300/r ), .b(\U1300/nback )
         );
    nand2_1 \U1300/U1103/U5  ( .x(\U1300/r ), .a(\U1300/naack ), .b(\U1300/s )
         );
    inv_1 \U1300/U1111/U3  ( .x(\U1300/reset ), .a(nbReset) );
    inv_1 \U1300/U1112/U3  ( .x(\U1300/naack ), .a(nba) );
    nor2_1 \U1300/U1130/U5  ( .x(\U1300/nback ), .a(nda), .b(\U1300/reset ) );
    aoai211_1 \U1300/U1128/U28/U1/U1  ( .x(\U1300/U1128/U28/U1/clr ), .a(
        \U1300/r ), .b(\U1300/naack ), .c(dg), .d(dsel) );
    nand3_1 \U1300/U1128/U28/U1/U2  ( .x(\U1300/U1128/U28/U1/set ), .a(dg), 
        .b(\U1300/r ), .c(\U1300/naack ) );
    nand2_2 \U1300/U1128/U28/U1/U3  ( .x(dsel), .a(\U1300/U1128/U28/U1/clr ), 
        .b(\U1300/U1128/U28/U1/set ) );
    aoai211_1 \U1300/U1127/U28/U1/U1  ( .x(\U1300/U1127/U28/U1/clr ), .a(
        \U1300/s ), .b(\U1300/nback ), .c(bg), .d(bsel) );
    nand3_1 \U1300/U1127/U28/U1/U2  ( .x(\U1300/U1127/U28/U1/set ), .a(bg), 
        .b(\U1300/s ), .c(\U1300/nback ) );
    nand2_2 \U1300/U1127/U28/U1/U3  ( .x(bsel), .a(\U1300/U1127/U28/U1/clr ), 
        .b(\U1300/U1127/U28/U1/set ) );
    aoai211_1 \U1289/U1150/U28/U1/U1  ( .x(\U1289/U1150/U28/U1/clr ), .a(il[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[2] ) );
    nand3_1 \U1289/U1150/U28/U1/U2  ( .x(\U1289/U1150/U28/U1/set ), .a(net195), 
        .b(il[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1150/U28/U1/U3  ( .x(\cdl[2] ), .a(
        \U1289/U1150/U28/U1/clr ), .b(\U1289/U1150/U28/U1/set ) );
    aoai211_1 \U1289/U1152/U28/U1/U1  ( .x(\U1289/U1152/U28/U1/clr ), .a(il[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[3] ) );
    nand3_1 \U1289/U1152/U28/U1/U2  ( .x(\U1289/U1152/U28/U1/set ), .a(net195), 
        .b(il[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1152/U28/U1/U3  ( .x(\cdl[3] ), .a(
        \U1289/U1152/U28/U1/clr ), .b(\U1289/U1152/U28/U1/set ) );
    aoai211_1 \U1289/U1149/U28/U1/U1  ( .x(\U1289/U1149/U28/U1/clr ), .a(ih[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[2] ) );
    nand3_1 \U1289/U1149/U28/U1/U2  ( .x(\U1289/U1149/U28/U1/set ), .a(net195), 
        .b(ih[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1149/U28/U1/U3  ( .x(\cdh[2] ), .a(
        \U1289/U1149/U28/U1/clr ), .b(\U1289/U1149/U28/U1/set ) );
    aoai211_1 \U1289/U1151/U28/U1/U1  ( .x(\U1289/U1151/U28/U1/clr ), .a(ih[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[3] ) );
    nand3_1 \U1289/U1151/U28/U1/U2  ( .x(\U1289/U1151/U28/U1/set ), .a(net195), 
        .b(ih[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1151/U28/U1/U3  ( .x(\cdh[3] ), .a(
        \U1289/U1151/U28/U1/clr ), .b(\U1289/U1151/U28/U1/set ) );
    inv_1 \U1289/U1148/U1147/U3  ( .x(\U1289/U1148/net189 ), .a(
        \U1289/bnreset ) );
    nor2_1 \U1289/U1148/U582/U5  ( .x(\U1289/U1148/net192 ), .a(\cdl[3] ), .b(
        \cdh[3] ) );
    nor2_1 \U1289/U1148/U580/U5  ( .x(\U1289/U1148/net191 ), .a(\cdl[2] ), .b(
        \cdh[2] ) );
    nor2_2 \U1289/U1148/U1146/U6  ( .x(\twobitack[2] ), .a(
        \U1289/U1148/net190 ), .b(\U1289/U1148/net189 ) );
    aoi222_1 \U1289/U1148/U1141/U30/U1  ( .x(\U1289/U1148/net190 ), .a(
        \U1289/U1148/net191 ), .b(\U1289/U1148/net192 ), .c(
        \U1289/U1148/net191 ), .d(\U1289/U1148/U1141/Z ), .e(
        \U1289/U1148/net192 ), .f(\U1289/U1148/U1141/Z ) );
    inv_1 \U1289/U1148/U1141/U30/Uinv  ( .x(\U1289/U1148/U1141/Z ), .a(
        \U1289/U1148/net190 ) );
    aoai211_1 \U1271/U1150/U28/U1/U1  ( .x(\U1271/U1150/U28/U1/clr ), .a(il[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[0] ) );
    nand3_1 \U1271/U1150/U28/U1/U2  ( .x(\U1271/U1150/U28/U1/set ), .a(net193), 
        .b(il[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1150/U28/U1/U3  ( .x(\cdl[0] ), .a(
        \U1271/U1150/U28/U1/clr ), .b(\U1271/U1150/U28/U1/set ) );
    aoai211_1 \U1271/U1152/U28/U1/U1  ( .x(\U1271/U1152/U28/U1/clr ), .a(il[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[1] ) );
    nand3_1 \U1271/U1152/U28/U1/U2  ( .x(\U1271/U1152/U28/U1/set ), .a(net193), 
        .b(il[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1152/U28/U1/U3  ( .x(\cdl[1] ), .a(
        \U1271/U1152/U28/U1/clr ), .b(\U1271/U1152/U28/U1/set ) );
    aoai211_1 \U1271/U1149/U28/U1/U1  ( .x(\U1271/U1149/U28/U1/clr ), .a(ih[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[0] ) );
    nand3_1 \U1271/U1149/U28/U1/U2  ( .x(\U1271/U1149/U28/U1/set ), .a(net193), 
        .b(ih[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1149/U28/U1/U3  ( .x(\cdh[0] ), .a(
        \U1271/U1149/U28/U1/clr ), .b(\U1271/U1149/U28/U1/set ) );
    aoai211_1 \U1271/U1151/U28/U1/U1  ( .x(\U1271/U1151/U28/U1/clr ), .a(ih[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[1] ) );
    nand3_1 \U1271/U1151/U28/U1/U2  ( .x(\U1271/U1151/U28/U1/set ), .a(net193), 
        .b(ih[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1151/U28/U1/U3  ( .x(\cdh[1] ), .a(
        \U1271/U1151/U28/U1/clr ), .b(\U1271/U1151/U28/U1/set ) );
    inv_1 \U1271/U1148/U1147/U3  ( .x(\U1271/U1148/net189 ), .a(
        \U1271/bnreset ) );
    nor2_1 \U1271/U1148/U582/U5  ( .x(\U1271/U1148/net192 ), .a(\cdl[1] ), .b(
        \cdh[1] ) );
    nor2_1 \U1271/U1148/U580/U5  ( .x(\U1271/U1148/net191 ), .a(\cdl[0] ), .b(
        \cdh[0] ) );
    nor2_2 \U1271/U1148/U1146/U6  ( .x(\twobitack[0] ), .a(
        \U1271/U1148/net190 ), .b(\U1271/U1148/net189 ) );
    aoi222_1 \U1271/U1148/U1141/U30/U1  ( .x(\U1271/U1148/net190 ), .a(
        \U1271/U1148/net191 ), .b(\U1271/U1148/net192 ), .c(
        \U1271/U1148/net191 ), .d(\U1271/U1148/U1141/Z ), .e(
        \U1271/U1148/net192 ), .f(\U1271/U1148/U1141/Z ) );
    inv_1 \U1271/U1148/U1141/U30/Uinv  ( .x(\U1271/U1148/U1141/Z ), .a(
        \U1271/U1148/net190 ) );
    nand2_1 \U1225/U1128/U5  ( .x(\U1225/s ), .a(\U1225/r ), .b(\U1225/nback )
         );
    nand2_1 \U1225/U1103/U5  ( .x(\U1225/r ), .a(\U1225/naack ), .b(\U1225/s )
         );
    inv_1 \U1225/U1111/U3  ( .x(\U1225/reset ), .a(nbReset) );
    inv_1 \U1225/U1112/U3  ( .x(\U1225/naack ), .a(nxa) );
    nor2_1 \U1225/U1127/U5  ( .x(\U1225/nback ), .a(nyla), .b(\U1225/reset )
         );
    and2_2 \U1225/U1129/U8  ( .x(xsel), .a(\U1225/nback ), .b(\U1225/s ) );
    and2_2 \U1225/U1124/U8  ( .x(ysel), .a(\U1225/r ), .b(\U1225/naack ) );
    and3_4 \U1308/U20/U9  ( .x(nya), .a(\U1308/nack[1] ), .b(\U1308/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U1308/U18/U5  ( .x(\U1308/nack[0] ), .a(\yl[3] ), .b(\yl[0] ) );
    nor2_1 \U1308/U19/U5  ( .x(\U1308/nack[1] ), .a(\yl[1] ), .b(\yl[2] ) );
    ao222_2 \U1308/U15_0_/U19/U1/U1  ( .x(\yl[0] ), .a(\y[0] ), .b(nyla), .c(
        \y[0] ), .d(\yl[0] ), .e(nyla), .f(\yl[0] ) );
    ao222_2 \U1308/U15_1_/U19/U1/U1  ( .x(\yl[1] ), .a(\y[1] ), .b(nyla), .c(
        \y[1] ), .d(\yl[1] ), .e(nyla), .f(\yl[1] ) );
    ao222_2 \U1308/U15_2_/U19/U1/U1  ( .x(\yl[2] ), .a(\y[2] ), .b(nyla), .c(
        \y[2] ), .d(\yl[2] ), .e(nyla), .f(\yl[2] ) );
    ao222_2 \U1308/U15_3_/U19/U1/U1  ( .x(\yl[3] ), .a(\y[3] ), .b(nyla), .c(
        \y[3] ), .d(\yl[3] ), .e(nyla), .f(\yl[3] ) );
    buf_3 U1 ( .x(\U1271/bnreset ), .a(nbReset) );
    buf_3 U2 ( .x(\U1289/bnreset ), .a(nbReset) );
endmodule


module chain_mergepackets_0 ( naa, nba, o, a, b, nReset, noa );
output [4:0] o;
input  [4:0] a;
input  [4:0] b;
input  nReset, noa;
output naa, nba;
    wire \noack[1] , \noack[0] , reset, bsel, as, setb, asel, seta, 
        \U916_0_/U25/U1/clr , \U916_0_/U25/U1/ob , \U916_1_/U25/U1/clr , 
        \U916_1_/U25/U1/ob , \U916_2_/U25/U1/clr , \U916_2_/U25/U1/ob , 
        \U916_3_/U25/U1/clr , \U916_3_/U25/U1/ob ;
    and2_1 \U1155/U8  ( .x(as), .a(seta), .b(asel) );
    nand2_1 \U1145/U5  ( .x(asel), .a(bsel), .b(seta) );
    nand2_1 \U1103/U5  ( .x(bsel), .a(setb), .b(asel) );
    inv_1 \U1135/U3  ( .x(reset), .a(nReset) );
    inv_1 \U1134/U3  ( .x(setb), .a(a[4]) );
    and3_2 \U1154/U9  ( .x(naa), .a(\noack[1] ), .b(\noack[0] ), .c(as) );
    nor3_1 \U1127/U7  ( .x(\noack[0] ), .a(o[1]), .b(reset), .c(o[0]) );
    nor2_1 \U1132/U5  ( .x(\noack[1] ), .a(o[3]), .b(o[2]) );
    oa31_1 \U916_0_/U25/U1/Uclr  ( .x(\U916_0_/U25/U1/clr ), .a(noa), .b(a[0]), 
        .c(b[0]), .d(o[0]) );
    oaoi211_1 \U916_0_/U25/U1/Uaoi  ( .x(\U916_0_/U25/U1/ob ), .a(a[0]), .b(b
        [0]), .c(noa), .d(\U916_0_/U25/U1/clr ) );
    inv_2 \U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U916_0_/U25/U1/ob ) );
    oa31_1 \U916_1_/U25/U1/Uclr  ( .x(\U916_1_/U25/U1/clr ), .a(noa), .b(a[1]), 
        .c(b[1]), .d(o[1]) );
    oaoi211_1 \U916_1_/U25/U1/Uaoi  ( .x(\U916_1_/U25/U1/ob ), .a(a[1]), .b(b
        [1]), .c(noa), .d(\U916_1_/U25/U1/clr ) );
    inv_2 \U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U916_1_/U25/U1/ob ) );
    oa31_1 \U916_2_/U25/U1/Uclr  ( .x(\U916_2_/U25/U1/clr ), .a(noa), .b(a[2]), 
        .c(b[2]), .d(o[2]) );
    oaoi211_1 \U916_2_/U25/U1/Uaoi  ( .x(\U916_2_/U25/U1/ob ), .a(a[2]), .b(b
        [2]), .c(noa), .d(\U916_2_/U25/U1/clr ) );
    inv_2 \U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U916_2_/U25/U1/ob ) );
    oa31_1 \U916_3_/U25/U1/Uclr  ( .x(\U916_3_/U25/U1/clr ), .a(noa), .b(a[3]), 
        .c(b[3]), .d(o[3]) );
    oaoi211_1 \U916_3_/U25/U1/Uaoi  ( .x(\U916_3_/U25/U1/ob ), .a(a[3]), .b(b
        [3]), .c(noa), .d(\U916_3_/U25/U1/clr ) );
    inv_2 \U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U916_3_/U25/U1/ob ) );
    ao222_2 \U1148/U19/U1/U1  ( .x(o[4]), .a(noa), .b(b[4]), .c(noa), .d(o[4]), 
        .e(b[4]), .f(o[4]) );
    aoi21_1 \U1153/U11  ( .x(seta), .a(o[4]), .b(setb), .c(reset) );
    and3_3 U1 ( .x(nba), .a(bsel), .b(\noack[0] ), .c(\noack[1] ) );
endmodule


module initiator_iport ( cack, chaincommand, err, nchainresponseack, nrouteack, 
    rd, routetxreq, rrnw, a, chainresponse, col, crnw, itag, lock, nReset, 
    nchaincommandack, pred, rack, route, routetxack, seq, size, wd );
output [4:0] chaincommand;
output [1:0] err;
output [63:0] rd;
output [1:0] rrnw;
input  [63:0] a;
input  [4:0] chainresponse;
input  [5:0] col;
input  [1:0] crnw;
input  [9:0] itag;
input  [1:0] lock;
input  [1:0] pred;
input  [4:0] route;
input  [1:0] seq;
input  [3:0] size;
input  [63:0] wd;
input  nReset, nchaincommandack, rack, routetxack;
output cack, nchainresponseack, nrouteack, routetxreq;
    wire \irbh[7] , \irbh[6] , \irbh[5] , \irbh[4] , \irbh[3] , \irbh[2] , 
        \irbh[1] , \irbh[0] , \ipayload[4] , \ipayload[3] , \ipayload[2] , 
        \ipayload[1] , \ipayload[0] , \icbh[7] , \icbh[6] , \icbh[5] , 
        \icbh[4] , \icbh[3] , \icbh[2] , \icbh[1] , \icbh[0] , \cstatus[1] , 
        \cstatus[0] , \irbl[7] , \irbl[6] , \irbl[5] , \irbl[4] , \irbl[3] , 
        \irbl[2] , \irbl[1] , \irbl[0] , \rstatus[1] , \rstatus[0] , 
        \can_defer[0] , \icbl[7] , \icbl[6] , \icbl[5] , \icbl[4] , \icbl[3] , 
        \icbl[2] , \icbl[1] , \icbl[0] , nircba, nResetb, responseack, 
        rstatusack, net165, reset, tok_ack, net170, ictrlack, icmdack, 
        ncstatusack, net116, pltxreq, net115, net128, pltxack, nicba, 
        nipayloadack, \U1662/U28/U1/clr , \U1662/U28/U1/set ;
    chain_irdemuxNew_0 U1442 ( .err(err), .ncback(nircba), .rd(rd), .rnw(rrnw), 
        .status({\rstatus[1] , \rstatus[0] }), .cbh({\irbh[7] , \irbh[6] , 
        \irbh[5] , \irbh[4] , \irbh[3] , \irbh[2] , \irbh[1] , \irbh[0] }), 
        .cbl({\irbl[7] , \irbl[6] , \irbl[5] , \irbl[4] , \irbl[3] , \irbl[2] , 
        \irbl[1] , \irbl[0] }), .nReset(nResetb), .nack(responseack), 
        .statusack(rstatusack) );
    chain_fr2dr_byte_3 chain_decoder ( .nia(nchainresponseack), .oh({\irbh[7] , 
        \irbh[6] , \irbh[5] , \irbh[4] , \irbh[3] , \irbh[2] , \irbh[1] , 
        \irbh[0] }), .ol({\irbl[7] , \irbl[6] , \irbl[5] , \irbl[4] , 
        \irbl[3] , \irbl[2] , \irbl[1] , \irbl[0] }), .i(chainresponse), 
        .nReset(nResetb), .noa(nircba) );
    chain_ic_ctrl_0 cmd_ctrl ( .ack(ictrlack), .candefer(\can_defer[0] ), 
        .eop(net116), .nstatack(ncstatusack), .pltxreq(pltxreq), .routetxreq(
        routetxreq), .tok_ack(tok_ack), .accept(\cstatus[0] ), .candefer_ack({
        1'b0, \can_defer[0] }), .defer(\cstatus[1] ), .eopack(net115), .lock(
        lock), .nReset(net128), .pltxack(pltxack), .routetxack(routetxack), 
        .tok_err(err[1]), .tok_ok(err[0]) );
    chain_icmux_0 cmd_mux ( .ack(icmdack), .chainh({\icbh[7] , \icbh[6] , 
        \icbh[5] , \icbh[4] , \icbh[3] , \icbh[2] , \icbh[1] , \icbh[0] }), 
        .chainl({\icbl[7] , \icbl[6] , \icbl[5] , \icbl[4] , \icbl[3] , 
        \icbl[2] , \icbl[1] , \icbl[0] }), .sendack(pltxack), .addr(a), .col(
        col), .itag(itag), .lock(lock), .nReset(net128), .nia(nicba), .pred(
        pred), .rnw(crnw), .sendreq(pltxreq), .seq(seq), .size(size), .wd(wd)
         );
    chain_dr2fr_byte_0 U1604 ( .eop_ack(net115), .ia(nicba), .o({\ipayload[4] , 
        \ipayload[3] , \ipayload[2] , \ipayload[1] , \ipayload[0] }), .eop(
        net116), .ih({\icbh[7] , \icbh[6] , \icbh[5] , \icbh[4] , \icbh[3] , 
        \icbh[2] , \icbh[1] , \icbh[0] }), .il({\icbl[7] , \icbl[6] , 
        \icbl[5] , \icbl[4] , \icbl[3] , \icbl[2] , \icbl[1] , \icbl[0] }), 
        .nReset(net128), .noa(nipayloadack) );
    chain_mergepackets_0 U1605 ( .naa(nrouteack), .nba(nipayloadack), .o(
        chaincommand), .a(route), .b({\ipayload[4] , \ipayload[3] , 
        \ipayload[2] , \ipayload[1] , \ipayload[0] }), .nReset(net128), .noa(
        nchaincommandack) );
    and2_1 U1676 ( .x(cack), .a(net170), .b(nResetb) );
    inv_4 \U1643/U3  ( .x(net128), .a(reset) );
    or2_4 \U1660/U12  ( .x(net165), .a(\cstatus[0] ), .b(\cstatus[1] ) );
    or2_1 \U1661/U12  ( .x(rstatusack), .a(net165), .b(reset) );
    ao222_2 \status_pipe_0_/U19/U1/U1  ( .x(\cstatus[0] ), .a(\rstatus[0] ), 
        .b(ncstatusack), .c(\rstatus[0] ), .d(\cstatus[0] ), .e(ncstatusack), 
        .f(\cstatus[0] ) );
    ao222_2 \status_pipe_1_/U19/U1/U1  ( .x(\cstatus[1] ), .a(\rstatus[1] ), 
        .b(ncstatusack), .c(\rstatus[1] ), .d(\cstatus[1] ), .e(ncstatusack), 
        .f(\cstatus[1] ) );
    ao222_1 \U1609/U18/U1/U1  ( .x(net170), .a(ictrlack), .b(icmdack), .c(
        ictrlack), .d(net170), .e(icmdack), .f(net170) );
    aoai211_1 \U1662/U28/U1/U1  ( .x(\U1662/U28/U1/clr ), .a(rack), .b(nResetb
        ), .c(tok_ack), .d(responseack) );
    nand3_1 \U1662/U28/U1/U2  ( .x(\U1662/U28/U1/set ), .a(tok_ack), .b(rack), 
        .c(nResetb) );
    nand2_2 \U1662/U28/U1/U3  ( .x(responseack), .a(\U1662/U28/U1/clr ), .b(
        \U1662/U28/U1/set ) );
    inv_2 U1 ( .x(reset), .a(nResetb) );
    buf_3 U2 ( .x(nResetb), .a(nReset) );
endmodule


module matched_delay_m2cp_com_iport ( x, a );
input  a;
output x;
    wire n2;
    buf_1 I1 ( .x(n2), .a(a) );
    buf_16 U1 ( .x(x), .a(n2) );
endmodule


module matched_delay_m2cp_resp_iport ( x, a );
input  a;
output x;
    assign x = a;
endmodule


module sr2dr_word_0 ( i, req, h, l );
input  [31:0] i;
output [31:0] h;
output [31:0] l;
input  req;
    wire \U31/nl , \U31/ni , \U31/nh , \U30/nl , \U30/ni , \U30/nh , \U29/nl , 
        \U29/ni , \U29/nh , \U28/nl , \U28/ni , \U28/nh , \U27/nl , \U27/ni , 
        \U27/nh , \U26/nl , \U26/ni , \U26/nh , \U25/nl , \U25/ni , \U25/nh , 
        \U24/nl , \U24/ni , \U24/nh , \U23/nl , \U23/ni , \U23/nh , \U22/nl , 
        \U22/ni , \U22/nh , \U21/nl , \U21/ni , \U21/nh , \U20/nl , \U20/ni , 
        \U20/nh , \U19/nl , \U19/ni , \U19/nh , \U18/nl , \U18/ni , \U18/nh , 
        \U17/nl , \U17/ni , \U17/nh , \U16/nl , \U16/ni , \U16/nh , \U15/nl , 
        \U15/ni , \U15/nh , \U14/nl , \U14/ni , \U14/nh , \U13/nl , \U13/ni , 
        \U13/nh , \U12/nl , \U12/ni , \U12/nh , \U11/nl , \U11/ni , \U11/nh , 
        \U10/nl , \U10/ni , \U10/nh , \U9/nl , \U9/ni , \U9/nh , \U8/nl , 
        \U8/ni , \U8/nh , \U7/nl , \U7/ni , \U7/nh , \U6/nl , \U6/ni , \U6/nh , 
        \U5/nl , \U5/ni , \U5/nh , \U4/nl , \U4/ni , \U4/nh , \U3/nl , \U3/ni , 
        \U3/nh , \U2/nl , \U2/ni , \U2/nh , \U1/nl , \U1/ni , \U1/nh , \U0/nl , 
        \U0/ni , \U0/nh , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
    inv_1 \U31/Uii  ( .x(\U31/ni ), .a(i[31]) );
    inv_1 \U31/Uih  ( .x(\U31/nh ), .a(h[31]) );
    inv_1 \U31/Uil  ( .x(\U31/nl ), .a(l[31]) );
    ao23_1 \U31/Ucl/U1/U1  ( .x(l[31]), .a(n9), .b(l[31]), .c(n1), .d(\U31/ni 
        ), .e(\U31/nh ) );
    ao23_1 \U31/Uch/U1/U1  ( .x(h[31]), .a(n9), .b(h[31]), .c(n2), .d(i[31]), 
        .e(\U31/nl ) );
    inv_1 \U30/Uii  ( .x(\U30/ni ), .a(i[30]) );
    inv_1 \U30/Uih  ( .x(\U30/nh ), .a(h[30]) );
    inv_1 \U30/Uil  ( .x(\U30/nl ), .a(l[30]) );
    ao23_1 \U30/Ucl/U1/U1  ( .x(l[30]), .a(n8), .b(l[30]), .c(n1), .d(\U30/ni 
        ), .e(\U30/nh ) );
    ao23_1 \U30/Uch/U1/U1  ( .x(h[30]), .a(n8), .b(h[30]), .c(n1), .d(i[30]), 
        .e(\U30/nl ) );
    inv_1 \U29/Uii  ( .x(\U29/ni ), .a(i[29]) );
    inv_1 \U29/Uih  ( .x(\U29/nh ), .a(h[29]) );
    inv_1 \U29/Uil  ( .x(\U29/nl ), .a(l[29]) );
    ao23_1 \U29/Ucl/U1/U1  ( .x(l[29]), .a(n8), .b(l[29]), .c(n1), .d(\U29/ni 
        ), .e(\U29/nh ) );
    ao23_1 \U29/Uch/U1/U1  ( .x(h[29]), .a(n8), .b(h[29]), .c(n2), .d(i[29]), 
        .e(\U29/nl ) );
    inv_1 \U28/Uii  ( .x(\U28/ni ), .a(i[28]) );
    inv_1 \U28/Uih  ( .x(\U28/nh ), .a(h[28]) );
    inv_1 \U28/Uil  ( .x(\U28/nl ), .a(l[28]) );
    ao23_1 \U28/Ucl/U1/U1  ( .x(l[28]), .a(n8), .b(l[28]), .c(n2), .d(\U28/ni 
        ), .e(\U28/nh ) );
    ao23_1 \U28/Uch/U1/U1  ( .x(h[28]), .a(n8), .b(h[28]), .c(n2), .d(i[28]), 
        .e(\U28/nl ) );
    inv_1 \U27/Uii  ( .x(\U27/ni ), .a(i[27]) );
    inv_1 \U27/Uih  ( .x(\U27/nh ), .a(h[27]) );
    inv_1 \U27/Uil  ( .x(\U27/nl ), .a(l[27]) );
    ao23_1 \U27/Ucl/U1/U1  ( .x(l[27]), .a(n8), .b(l[27]), .c(n2), .d(\U27/ni 
        ), .e(\U27/nh ) );
    ao23_1 \U27/Uch/U1/U1  ( .x(h[27]), .a(n8), .b(h[27]), .c(n2), .d(i[27]), 
        .e(\U27/nl ) );
    inv_1 \U26/Uii  ( .x(\U26/ni ), .a(i[26]) );
    inv_1 \U26/Uih  ( .x(\U26/nh ), .a(h[26]) );
    inv_1 \U26/Uil  ( .x(\U26/nl ), .a(l[26]) );
    ao23_1 \U26/Ucl/U1/U1  ( .x(l[26]), .a(n7), .b(l[26]), .c(n2), .d(\U26/ni 
        ), .e(\U26/nh ) );
    ao23_1 \U26/Uch/U1/U1  ( .x(h[26]), .a(n7), .b(h[26]), .c(n4), .d(i[26]), 
        .e(\U26/nl ) );
    inv_1 \U25/Uii  ( .x(\U25/ni ), .a(i[25]) );
    inv_1 \U25/Uih  ( .x(\U25/nh ), .a(h[25]) );
    inv_1 \U25/Uil  ( .x(\U25/nl ), .a(l[25]) );
    ao23_1 \U25/Ucl/U1/U1  ( .x(l[25]), .a(n7), .b(l[25]), .c(n4), .d(\U25/ni 
        ), .e(\U25/nh ) );
    ao23_1 \U25/Uch/U1/U1  ( .x(h[25]), .a(n7), .b(h[25]), .c(n4), .d(i[25]), 
        .e(\U25/nl ) );
    inv_1 \U24/Uii  ( .x(\U24/ni ), .a(i[24]) );
    inv_1 \U24/Uih  ( .x(\U24/nh ), .a(h[24]) );
    inv_1 \U24/Uil  ( .x(\U24/nl ), .a(l[24]) );
    ao23_1 \U24/Ucl/U1/U1  ( .x(l[24]), .a(n7), .b(l[24]), .c(n4), .d(\U24/ni 
        ), .e(\U24/nh ) );
    ao23_1 \U24/Uch/U1/U1  ( .x(h[24]), .a(n7), .b(h[24]), .c(n4), .d(i[24]), 
        .e(\U24/nl ) );
    inv_1 \U23/Uii  ( .x(\U23/ni ), .a(i[23]) );
    inv_1 \U23/Uih  ( .x(\U23/nh ), .a(h[23]) );
    inv_1 \U23/Uil  ( .x(\U23/nl ), .a(l[23]) );
    ao23_1 \U23/Ucl/U1/U1  ( .x(l[23]), .a(n7), .b(l[23]), .c(n3), .d(\U23/ni 
        ), .e(\U23/nh ) );
    ao23_1 \U23/Uch/U1/U1  ( .x(h[23]), .a(n7), .b(h[23]), .c(n3), .d(i[23]), 
        .e(\U23/nl ) );
    inv_1 \U22/Uii  ( .x(\U22/ni ), .a(i[22]) );
    inv_1 \U22/Uih  ( .x(\U22/nh ), .a(h[22]) );
    inv_1 \U22/Uil  ( .x(\U22/nl ), .a(l[22]) );
    ao23_1 \U22/Ucl/U1/U1  ( .x(l[22]), .a(n6), .b(l[22]), .c(n3), .d(\U22/ni 
        ), .e(\U22/nh ) );
    ao23_1 \U22/Uch/U1/U1  ( .x(h[22]), .a(n6), .b(h[22]), .c(n3), .d(i[22]), 
        .e(\U22/nl ) );
    inv_1 \U21/Uii  ( .x(\U21/ni ), .a(i[21]) );
    inv_1 \U21/Uih  ( .x(\U21/nh ), .a(h[21]) );
    inv_1 \U21/Uil  ( .x(\U21/nl ), .a(l[21]) );
    ao23_1 \U21/Ucl/U1/U1  ( .x(l[21]), .a(n6), .b(l[21]), .c(n3), .d(\U21/ni 
        ), .e(\U21/nh ) );
    ao23_1 \U21/Uch/U1/U1  ( .x(h[21]), .a(n6), .b(h[21]), .c(n3), .d(i[21]), 
        .e(\U21/nl ) );
    inv_1 \U20/Uii  ( .x(\U20/ni ), .a(i[20]) );
    inv_1 \U20/Uih  ( .x(\U20/nh ), .a(h[20]) );
    inv_1 \U20/Uil  ( .x(\U20/nl ), .a(l[20]) );
    ao23_1 \U20/Ucl/U1/U1  ( .x(l[20]), .a(n6), .b(l[20]), .c(n5), .d(\U20/ni 
        ), .e(\U20/nh ) );
    ao23_1 \U20/Uch/U1/U1  ( .x(h[20]), .a(n6), .b(h[20]), .c(n4), .d(i[20]), 
        .e(\U20/nl ) );
    inv_1 \U19/Uii  ( .x(\U19/ni ), .a(i[19]) );
    inv_1 \U19/Uih  ( .x(\U19/nh ), .a(h[19]) );
    inv_1 \U19/Uil  ( .x(\U19/nl ), .a(l[19]) );
    ao23_1 \U19/Ucl/U1/U1  ( .x(l[19]), .a(n6), .b(l[19]), .c(n4), .d(\U19/ni 
        ), .e(\U19/nh ) );
    ao23_1 \U19/Uch/U1/U1  ( .x(h[19]), .a(n6), .b(h[19]), .c(n4), .d(i[19]), 
        .e(\U19/nl ) );
    inv_1 \U18/Uii  ( .x(\U18/ni ), .a(i[18]) );
    inv_1 \U18/Uih  ( .x(\U18/nh ), .a(h[18]) );
    inv_1 \U18/Uil  ( .x(\U18/nl ), .a(l[18]) );
    ao23_1 \U18/Ucl/U1/U1  ( .x(l[18]), .a(n5), .b(l[18]), .c(n5), .d(\U18/ni 
        ), .e(\U18/nh ) );
    ao23_1 \U18/Uch/U1/U1  ( .x(h[18]), .a(n5), .b(h[18]), .c(n5), .d(i[18]), 
        .e(\U18/nl ) );
    inv_1 \U17/Uii  ( .x(\U17/ni ), .a(i[17]) );
    inv_1 \U17/Uih  ( .x(\U17/nh ), .a(h[17]) );
    inv_1 \U17/Uil  ( .x(\U17/nl ), .a(l[17]) );
    ao23_1 \U17/Ucl/U1/U1  ( .x(l[17]), .a(n6), .b(l[17]), .c(n5), .d(\U17/ni 
        ), .e(\U17/nh ) );
    ao23_1 \U17/Uch/U1/U1  ( .x(h[17]), .a(n7), .b(h[17]), .c(n4), .d(i[17]), 
        .e(\U17/nl ) );
    inv_1 \U16/Uii  ( .x(\U16/ni ), .a(i[16]) );
    inv_1 \U16/Uih  ( .x(\U16/nh ), .a(h[16]) );
    inv_1 \U16/Uil  ( .x(\U16/nl ), .a(l[16]) );
    ao23_1 \U16/Ucl/U1/U1  ( .x(l[16]), .a(n9), .b(l[16]), .c(n3), .d(\U16/ni 
        ), .e(\U16/nh ) );
    ao23_1 \U16/Uch/U1/U1  ( .x(h[16]), .a(n9), .b(h[16]), .c(n1), .d(i[16]), 
        .e(\U16/nl ) );
    inv_1 \U15/Uii  ( .x(\U15/ni ), .a(i[15]) );
    inv_1 \U15/Uih  ( .x(\U15/nh ), .a(h[15]) );
    inv_1 \U15/Uil  ( .x(\U15/nl ), .a(l[15]) );
    ao23_1 \U15/Ucl/U1/U1  ( .x(l[15]), .a(n8), .b(l[15]), .c(n1), .d(\U15/ni 
        ), .e(\U15/nh ) );
    ao23_1 \U15/Uch/U1/U1  ( .x(h[15]), .a(n7), .b(h[15]), .c(n1), .d(i[15]), 
        .e(\U15/nl ) );
    inv_1 \U14/Uii  ( .x(\U14/ni ), .a(i[14]) );
    inv_1 \U14/Uih  ( .x(\U14/nh ), .a(h[14]) );
    inv_1 \U14/Uil  ( .x(\U14/nl ), .a(l[14]) );
    ao23_1 \U14/Ucl/U1/U1  ( .x(l[14]), .a(n6), .b(l[14]), .c(n1), .d(\U14/ni 
        ), .e(\U14/nh ) );
    ao23_1 \U14/Uch/U1/U1  ( .x(h[14]), .a(n6), .b(h[14]), .c(n3), .d(i[14]), 
        .e(\U14/nl ) );
    inv_1 \U13/Uii  ( .x(\U13/ni ), .a(i[13]) );
    inv_1 \U13/Uih  ( .x(\U13/nh ), .a(h[13]) );
    inv_1 \U13/Uil  ( .x(\U13/nl ), .a(l[13]) );
    ao23_1 \U13/Ucl/U1/U1  ( .x(l[13]), .a(n6), .b(l[13]), .c(n4), .d(\U13/ni 
        ), .e(\U13/nh ) );
    ao23_1 \U13/Uch/U1/U1  ( .x(h[13]), .a(n6), .b(h[13]), .c(n4), .d(i[13]), 
        .e(\U13/nl ) );
    inv_1 \U12/Uii  ( .x(\U12/ni ), .a(i[12]) );
    inv_1 \U12/Uih  ( .x(\U12/nh ), .a(h[12]) );
    inv_1 \U12/Uil  ( .x(\U12/nl ), .a(l[12]) );
    ao23_1 \U12/Ucl/U1/U1  ( .x(l[12]), .a(n5), .b(l[12]), .c(n4), .d(\U12/ni 
        ), .e(\U12/nh ) );
    ao23_1 \U12/Uch/U1/U1  ( .x(h[12]), .a(n5), .b(h[12]), .c(n4), .d(i[12]), 
        .e(\U12/nl ) );
    inv_1 \U11/Uii  ( .x(\U11/ni ), .a(i[11]) );
    inv_1 \U11/Uih  ( .x(\U11/nh ), .a(h[11]) );
    inv_1 \U11/Uil  ( .x(\U11/nl ), .a(l[11]) );
    ao23_1 \U11/Ucl/U1/U1  ( .x(l[11]), .a(n5), .b(l[11]), .c(n4), .d(\U11/ni 
        ), .e(\U11/nh ) );
    ao23_1 \U11/Uch/U1/U1  ( .x(h[11]), .a(n5), .b(h[11]), .c(n4), .d(i[11]), 
        .e(\U11/nl ) );
    inv_1 \U10/Uii  ( .x(\U10/ni ), .a(i[10]) );
    inv_1 \U10/Uih  ( .x(\U10/nh ), .a(h[10]) );
    inv_1 \U10/Uil  ( .x(\U10/nl ), .a(l[10]) );
    ao23_1 \U10/Ucl/U1/U1  ( .x(l[10]), .a(n5), .b(l[10]), .c(n3), .d(\U10/ni 
        ), .e(\U10/nh ) );
    ao23_1 \U10/Uch/U1/U1  ( .x(h[10]), .a(n5), .b(h[10]), .c(n3), .d(i[10]), 
        .e(\U10/nl ) );
    inv_1 \U9/Uii  ( .x(\U9/ni ), .a(i[9]) );
    inv_1 \U9/Uih  ( .x(\U9/nh ), .a(h[9]) );
    inv_1 \U9/Uil  ( .x(\U9/nl ), .a(l[9]) );
    ao23_1 \U9/Ucl/U1/U1  ( .x(l[9]), .a(n5), .b(l[9]), .c(n3), .d(\U9/ni ), 
        .e(\U9/nh ) );
    ao23_1 \U9/Uch/U1/U1  ( .x(h[9]), .a(n5), .b(h[9]), .c(n3), .d(i[9]), .e(
        \U9/nl ) );
    inv_1 \U8/Uii  ( .x(\U8/ni ), .a(i[8]) );
    inv_1 \U8/Uih  ( .x(\U8/nh ), .a(h[8]) );
    inv_1 \U8/Uil  ( .x(\U8/nl ), .a(l[8]) );
    ao23_1 \U8/Ucl/U1/U1  ( .x(l[8]), .a(n5), .b(l[8]), .c(n3), .d(\U8/ni ), 
        .e(\U8/nh ) );
    ao23_1 \U8/Uch/U1/U1  ( .x(h[8]), .a(n5), .b(h[8]), .c(n3), .d(i[8]), .e(
        \U8/nl ) );
    inv_1 \U7/Uii  ( .x(\U7/ni ), .a(i[7]) );
    inv_1 \U7/Uih  ( .x(\U7/nh ), .a(h[7]) );
    inv_1 \U7/Uil  ( .x(\U7/nl ), .a(l[7]) );
    ao23_1 \U7/Ucl/U1/U1  ( .x(l[7]), .a(n7), .b(l[7]), .c(n3), .d(\U7/ni ), 
        .e(\U7/nh ) );
    ao23_1 \U7/Uch/U1/U1  ( .x(h[7]), .a(n7), .b(h[7]), .c(n2), .d(i[7]), .e(
        \U7/nl ) );
    inv_1 \U6/Uii  ( .x(\U6/ni ), .a(i[6]) );
    inv_1 \U6/Uih  ( .x(\U6/nh ), .a(h[6]) );
    inv_1 \U6/Uil  ( .x(\U6/nl ), .a(l[6]) );
    ao23_1 \U6/Ucl/U1/U1  ( .x(l[6]), .a(n7), .b(l[6]), .c(n2), .d(\U6/ni ), 
        .e(\U6/nh ) );
    ao23_1 \U6/Uch/U1/U1  ( .x(h[6]), .a(n7), .b(h[6]), .c(n2), .d(i[6]), .e(
        \U6/nl ) );
    inv_1 \U5/Uii  ( .x(\U5/ni ), .a(i[5]) );
    inv_1 \U5/Uih  ( .x(\U5/nh ), .a(h[5]) );
    inv_1 \U5/Uil  ( .x(\U5/nl ), .a(l[5]) );
    ao23_1 \U5/Ucl/U1/U1  ( .x(l[5]), .a(n7), .b(l[5]), .c(n2), .d(\U5/ni ), 
        .e(\U5/nh ) );
    ao23_1 \U5/Uch/U1/U1  ( .x(h[5]), .a(n7), .b(h[5]), .c(n2), .d(i[5]), .e(
        \U5/nl ) );
    inv_1 \U4/Uii  ( .x(\U4/ni ), .a(i[4]) );
    inv_1 \U4/Uih  ( .x(\U4/nh ), .a(h[4]) );
    inv_1 \U4/Uil  ( .x(\U4/nl ), .a(l[4]) );
    ao23_1 \U4/Ucl/U1/U1  ( .x(l[4]), .a(n6), .b(l[4]), .c(n2), .d(\U4/ni ), 
        .e(\U4/nh ) );
    ao23_1 \U4/Uch/U1/U1  ( .x(h[4]), .a(n6), .b(h[4]), .c(n2), .d(i[4]), .e(
        \U4/nl ) );
    inv_1 \U3/Uii  ( .x(\U3/ni ), .a(i[3]) );
    inv_1 \U3/Uih  ( .x(\U3/nh ), .a(h[3]) );
    inv_1 \U3/Uil  ( .x(\U3/nl ), .a(l[3]) );
    ao23_1 \U3/Ucl/U1/U1  ( .x(l[3]), .a(n6), .b(l[3]), .c(n2), .d(\U3/ni ), 
        .e(\U3/nh ) );
    ao23_1 \U3/Uch/U1/U1  ( .x(h[3]), .a(n8), .b(h[3]), .c(n1), .d(i[3]), .e(
        \U3/nl ) );
    inv_1 \U2/Uii  ( .x(\U2/ni ), .a(i[2]) );
    inv_1 \U2/Uih  ( .x(\U2/nh ), .a(h[2]) );
    inv_1 \U2/Uil  ( .x(\U2/nl ), .a(l[2]) );
    ao23_1 \U2/Ucl/U1/U1  ( .x(l[2]), .a(n8), .b(l[2]), .c(n1), .d(\U2/ni ), 
        .e(\U2/nh ) );
    ao23_1 \U2/Uch/U1/U1  ( .x(h[2]), .a(n8), .b(h[2]), .c(n1), .d(i[2]), .e(
        \U2/nl ) );
    inv_1 \U1/Uii  ( .x(\U1/ni ), .a(i[1]) );
    inv_1 \U1/Uih  ( .x(\U1/nh ), .a(h[1]) );
    inv_1 \U1/Uil  ( .x(\U1/nl ), .a(l[1]) );
    ao23_1 \U1/Ucl/U1/U1  ( .x(l[1]), .a(n8), .b(l[1]), .c(n1), .d(\U1/ni ), 
        .e(\U1/nh ) );
    ao23_1 \U1/Uch/U1/U1  ( .x(h[1]), .a(n8), .b(h[1]), .c(n1), .d(i[1]), .e(
        \U1/nl ) );
    inv_1 \U0/Uii  ( .x(\U0/ni ), .a(i[0]) );
    inv_1 \U0/Uih  ( .x(\U0/nh ), .a(h[0]) );
    inv_1 \U0/Uil  ( .x(\U0/nl ), .a(l[0]) );
    ao23_1 \U0/Ucl/U1/U1  ( .x(l[0]), .a(n8), .b(l[0]), .c(n1), .d(\U0/ni ), 
        .e(\U0/nh ) );
    ao23_1 \U0/Uch/U1/U1  ( .x(h[0]), .a(n8), .b(h[0]), .c(n1), .d(i[0]), .e(
        \U0/nl ) );
    buf_16 U1 ( .x(n1), .a(n12) );
    buf_16 U2 ( .x(n2), .a(n12) );
    buf_16 U3 ( .x(n3), .a(n12) );
    buf_16 U4 ( .x(n4), .a(n11) );
    buf_16 U5 ( .x(n5), .a(n11) );
    buf_16 U6 ( .x(n6), .a(n11) );
    buf_16 U7 ( .x(n7), .a(n10) );
    buf_16 U8 ( .x(n8), .a(n10) );
    buf_16 U9 ( .x(n9), .a(n10) );
    buf_16 U10 ( .x(n10), .a(req) );
    buf_16 U11 ( .x(n11), .a(req) );
    buf_16 U12 ( .x(n12), .a(req) );
endmodule


module sr2dr_word_1 ( i, req, h, l );
input  [31:0] i;
output [31:0] h;
output [31:0] l;
input  req;
    wire \U31/nl , \U31/ni , \U31/nh , \U30/nl , \U30/ni , \U30/nh , \U29/nl , 
        \U29/ni , \U29/nh , \U28/nl , \U28/ni , \U28/nh , \U27/nl , \U27/ni , 
        \U27/nh , \U26/nl , \U26/ni , \U26/nh , \U25/nl , \U25/ni , \U25/nh , 
        \U24/nl , \U24/ni , \U24/nh , \U23/nl , \U23/ni , \U23/nh , \U22/nl , 
        \U22/ni , \U22/nh , \U21/nl , \U21/ni , \U21/nh , \U20/nl , \U20/ni , 
        \U20/nh , \U19/nl , \U19/ni , \U19/nh , \U18/nl , \U18/ni , \U18/nh , 
        \U17/nl , \U17/ni , \U17/nh , \U16/nl , \U16/ni , \U16/nh , \U15/nl , 
        \U15/ni , \U15/nh , \U14/nl , \U14/ni , \U14/nh , \U13/nl , \U13/ni , 
        \U13/nh , \U12/nl , \U12/ni , \U12/nh , \U11/nl , \U11/ni , \U11/nh , 
        \U10/nl , \U10/ni , \U10/nh , \U9/nl , \U9/ni , \U9/nh , \U8/nl , 
        \U8/ni , \U8/nh , \U7/nl , \U7/ni , \U7/nh , \U6/nl , \U6/ni , \U6/nh , 
        \U5/nl , \U5/ni , \U5/nh , \U4/nl , \U4/ni , \U4/nh , \U3/nl , \U3/ni , 
        \U3/nh , \U2/nl , \U2/ni , \U2/nh , \U1/nl , \U1/ni , \U1/nh , \U0/nl , 
        \U0/ni , \U0/nh , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
    inv_1 \U31/Uii  ( .x(\U31/ni ), .a(i[31]) );
    inv_1 \U31/Uih  ( .x(\U31/nh ), .a(h[31]) );
    inv_1 \U31/Uil  ( .x(\U31/nl ), .a(l[31]) );
    ao23_1 \U31/Ucl/U1/U1  ( .x(l[31]), .a(n9), .b(l[31]), .c(n1), .d(\U31/ni 
        ), .e(\U31/nh ) );
    ao23_1 \U31/Uch/U1/U1  ( .x(h[31]), .a(n9), .b(h[31]), .c(n2), .d(i[31]), 
        .e(\U31/nl ) );
    inv_1 \U30/Uii  ( .x(\U30/ni ), .a(i[30]) );
    inv_1 \U30/Uih  ( .x(\U30/nh ), .a(h[30]) );
    inv_1 \U30/Uil  ( .x(\U30/nl ), .a(l[30]) );
    ao23_1 \U30/Ucl/U1/U1  ( .x(l[30]), .a(n8), .b(l[30]), .c(n1), .d(\U30/ni 
        ), .e(\U30/nh ) );
    ao23_1 \U30/Uch/U1/U1  ( .x(h[30]), .a(n8), .b(h[30]), .c(n1), .d(i[30]), 
        .e(\U30/nl ) );
    inv_1 \U29/Uii  ( .x(\U29/ni ), .a(i[29]) );
    inv_1 \U29/Uih  ( .x(\U29/nh ), .a(h[29]) );
    inv_1 \U29/Uil  ( .x(\U29/nl ), .a(l[29]) );
    ao23_1 \U29/Ucl/U1/U1  ( .x(l[29]), .a(n8), .b(l[29]), .c(n1), .d(\U29/ni 
        ), .e(\U29/nh ) );
    ao23_1 \U29/Uch/U1/U1  ( .x(h[29]), .a(n8), .b(h[29]), .c(n2), .d(i[29]), 
        .e(\U29/nl ) );
    inv_1 \U28/Uii  ( .x(\U28/ni ), .a(i[28]) );
    inv_1 \U28/Uih  ( .x(\U28/nh ), .a(h[28]) );
    inv_1 \U28/Uil  ( .x(\U28/nl ), .a(l[28]) );
    ao23_1 \U28/Ucl/U1/U1  ( .x(l[28]), .a(n8), .b(l[28]), .c(n2), .d(\U28/ni 
        ), .e(\U28/nh ) );
    ao23_1 \U28/Uch/U1/U1  ( .x(h[28]), .a(n8), .b(h[28]), .c(n2), .d(i[28]), 
        .e(\U28/nl ) );
    inv_1 \U27/Uii  ( .x(\U27/ni ), .a(i[27]) );
    inv_1 \U27/Uih  ( .x(\U27/nh ), .a(h[27]) );
    inv_1 \U27/Uil  ( .x(\U27/nl ), .a(l[27]) );
    ao23_1 \U27/Ucl/U1/U1  ( .x(l[27]), .a(n8), .b(l[27]), .c(n2), .d(\U27/ni 
        ), .e(\U27/nh ) );
    ao23_1 \U27/Uch/U1/U1  ( .x(h[27]), .a(n8), .b(h[27]), .c(n2), .d(i[27]), 
        .e(\U27/nl ) );
    inv_1 \U26/Uii  ( .x(\U26/ni ), .a(i[26]) );
    inv_1 \U26/Uih  ( .x(\U26/nh ), .a(h[26]) );
    inv_1 \U26/Uil  ( .x(\U26/nl ), .a(l[26]) );
    ao23_1 \U26/Ucl/U1/U1  ( .x(l[26]), .a(n7), .b(l[26]), .c(n2), .d(\U26/ni 
        ), .e(\U26/nh ) );
    ao23_1 \U26/Uch/U1/U1  ( .x(h[26]), .a(n7), .b(h[26]), .c(n4), .d(i[26]), 
        .e(\U26/nl ) );
    inv_1 \U25/Uii  ( .x(\U25/ni ), .a(i[25]) );
    inv_1 \U25/Uih  ( .x(\U25/nh ), .a(h[25]) );
    inv_1 \U25/Uil  ( .x(\U25/nl ), .a(l[25]) );
    ao23_1 \U25/Ucl/U1/U1  ( .x(l[25]), .a(n7), .b(l[25]), .c(n4), .d(\U25/ni 
        ), .e(\U25/nh ) );
    ao23_1 \U25/Uch/U1/U1  ( .x(h[25]), .a(n7), .b(h[25]), .c(n4), .d(i[25]), 
        .e(\U25/nl ) );
    inv_1 \U24/Uii  ( .x(\U24/ni ), .a(i[24]) );
    inv_1 \U24/Uih  ( .x(\U24/nh ), .a(h[24]) );
    inv_1 \U24/Uil  ( .x(\U24/nl ), .a(l[24]) );
    ao23_1 \U24/Ucl/U1/U1  ( .x(l[24]), .a(n7), .b(l[24]), .c(n4), .d(\U24/ni 
        ), .e(\U24/nh ) );
    ao23_1 \U24/Uch/U1/U1  ( .x(h[24]), .a(n7), .b(h[24]), .c(n4), .d(i[24]), 
        .e(\U24/nl ) );
    inv_1 \U23/Uii  ( .x(\U23/ni ), .a(i[23]) );
    inv_1 \U23/Uih  ( .x(\U23/nh ), .a(h[23]) );
    inv_1 \U23/Uil  ( .x(\U23/nl ), .a(l[23]) );
    ao23_1 \U23/Ucl/U1/U1  ( .x(l[23]), .a(n7), .b(l[23]), .c(n3), .d(\U23/ni 
        ), .e(\U23/nh ) );
    ao23_1 \U23/Uch/U1/U1  ( .x(h[23]), .a(n7), .b(h[23]), .c(n3), .d(i[23]), 
        .e(\U23/nl ) );
    inv_1 \U22/Uii  ( .x(\U22/ni ), .a(i[22]) );
    inv_1 \U22/Uih  ( .x(\U22/nh ), .a(h[22]) );
    inv_1 \U22/Uil  ( .x(\U22/nl ), .a(l[22]) );
    ao23_1 \U22/Ucl/U1/U1  ( .x(l[22]), .a(n6), .b(l[22]), .c(n3), .d(\U22/ni 
        ), .e(\U22/nh ) );
    ao23_1 \U22/Uch/U1/U1  ( .x(h[22]), .a(n6), .b(h[22]), .c(n3), .d(i[22]), 
        .e(\U22/nl ) );
    inv_1 \U21/Uii  ( .x(\U21/ni ), .a(i[21]) );
    inv_1 \U21/Uih  ( .x(\U21/nh ), .a(h[21]) );
    inv_1 \U21/Uil  ( .x(\U21/nl ), .a(l[21]) );
    ao23_1 \U21/Ucl/U1/U1  ( .x(l[21]), .a(n6), .b(l[21]), .c(n3), .d(\U21/ni 
        ), .e(\U21/nh ) );
    ao23_1 \U21/Uch/U1/U1  ( .x(h[21]), .a(n6), .b(h[21]), .c(n3), .d(i[21]), 
        .e(\U21/nl ) );
    inv_1 \U20/Uii  ( .x(\U20/ni ), .a(i[20]) );
    inv_1 \U20/Uih  ( .x(\U20/nh ), .a(h[20]) );
    inv_1 \U20/Uil  ( .x(\U20/nl ), .a(l[20]) );
    ao23_1 \U20/Ucl/U1/U1  ( .x(l[20]), .a(n6), .b(l[20]), .c(n5), .d(\U20/ni 
        ), .e(\U20/nh ) );
    ao23_1 \U20/Uch/U1/U1  ( .x(h[20]), .a(n6), .b(h[20]), .c(n4), .d(i[20]), 
        .e(\U20/nl ) );
    inv_1 \U19/Uii  ( .x(\U19/ni ), .a(i[19]) );
    inv_1 \U19/Uih  ( .x(\U19/nh ), .a(h[19]) );
    inv_1 \U19/Uil  ( .x(\U19/nl ), .a(l[19]) );
    ao23_1 \U19/Ucl/U1/U1  ( .x(l[19]), .a(n6), .b(l[19]), .c(n4), .d(\U19/ni 
        ), .e(\U19/nh ) );
    ao23_1 \U19/Uch/U1/U1  ( .x(h[19]), .a(n6), .b(h[19]), .c(n4), .d(i[19]), 
        .e(\U19/nl ) );
    inv_1 \U18/Uii  ( .x(\U18/ni ), .a(i[18]) );
    inv_1 \U18/Uih  ( .x(\U18/nh ), .a(h[18]) );
    inv_1 \U18/Uil  ( .x(\U18/nl ), .a(l[18]) );
    ao23_1 \U18/Ucl/U1/U1  ( .x(l[18]), .a(n5), .b(l[18]), .c(n5), .d(\U18/ni 
        ), .e(\U18/nh ) );
    ao23_1 \U18/Uch/U1/U1  ( .x(h[18]), .a(n5), .b(h[18]), .c(n5), .d(i[18]), 
        .e(\U18/nl ) );
    inv_1 \U17/Uii  ( .x(\U17/ni ), .a(i[17]) );
    inv_1 \U17/Uih  ( .x(\U17/nh ), .a(h[17]) );
    inv_1 \U17/Uil  ( .x(\U17/nl ), .a(l[17]) );
    ao23_1 \U17/Ucl/U1/U1  ( .x(l[17]), .a(n6), .b(l[17]), .c(n5), .d(\U17/ni 
        ), .e(\U17/nh ) );
    ao23_1 \U17/Uch/U1/U1  ( .x(h[17]), .a(n7), .b(h[17]), .c(n4), .d(i[17]), 
        .e(\U17/nl ) );
    inv_1 \U16/Uii  ( .x(\U16/ni ), .a(i[16]) );
    inv_1 \U16/Uih  ( .x(\U16/nh ), .a(h[16]) );
    inv_1 \U16/Uil  ( .x(\U16/nl ), .a(l[16]) );
    ao23_1 \U16/Ucl/U1/U1  ( .x(l[16]), .a(n9), .b(l[16]), .c(n3), .d(\U16/ni 
        ), .e(\U16/nh ) );
    ao23_1 \U16/Uch/U1/U1  ( .x(h[16]), .a(n9), .b(h[16]), .c(n1), .d(i[16]), 
        .e(\U16/nl ) );
    inv_1 \U15/Uii  ( .x(\U15/ni ), .a(i[15]) );
    inv_1 \U15/Uih  ( .x(\U15/nh ), .a(h[15]) );
    inv_1 \U15/Uil  ( .x(\U15/nl ), .a(l[15]) );
    ao23_1 \U15/Ucl/U1/U1  ( .x(l[15]), .a(n8), .b(l[15]), .c(n1), .d(\U15/ni 
        ), .e(\U15/nh ) );
    ao23_1 \U15/Uch/U1/U1  ( .x(h[15]), .a(n7), .b(h[15]), .c(n1), .d(i[15]), 
        .e(\U15/nl ) );
    inv_1 \U14/Uii  ( .x(\U14/ni ), .a(i[14]) );
    inv_1 \U14/Uih  ( .x(\U14/nh ), .a(h[14]) );
    inv_1 \U14/Uil  ( .x(\U14/nl ), .a(l[14]) );
    ao23_1 \U14/Ucl/U1/U1  ( .x(l[14]), .a(n6), .b(l[14]), .c(n1), .d(\U14/ni 
        ), .e(\U14/nh ) );
    ao23_1 \U14/Uch/U1/U1  ( .x(h[14]), .a(n6), .b(h[14]), .c(n3), .d(i[14]), 
        .e(\U14/nl ) );
    inv_1 \U13/Uii  ( .x(\U13/ni ), .a(i[13]) );
    inv_1 \U13/Uih  ( .x(\U13/nh ), .a(h[13]) );
    inv_1 \U13/Uil  ( .x(\U13/nl ), .a(l[13]) );
    ao23_1 \U13/Ucl/U1/U1  ( .x(l[13]), .a(n6), .b(l[13]), .c(n4), .d(\U13/ni 
        ), .e(\U13/nh ) );
    ao23_1 \U13/Uch/U1/U1  ( .x(h[13]), .a(n6), .b(h[13]), .c(n4), .d(i[13]), 
        .e(\U13/nl ) );
    inv_1 \U12/Uii  ( .x(\U12/ni ), .a(i[12]) );
    inv_1 \U12/Uih  ( .x(\U12/nh ), .a(h[12]) );
    inv_1 \U12/Uil  ( .x(\U12/nl ), .a(l[12]) );
    ao23_1 \U12/Ucl/U1/U1  ( .x(l[12]), .a(n5), .b(l[12]), .c(n4), .d(\U12/ni 
        ), .e(\U12/nh ) );
    ao23_1 \U12/Uch/U1/U1  ( .x(h[12]), .a(n5), .b(h[12]), .c(n4), .d(i[12]), 
        .e(\U12/nl ) );
    inv_1 \U11/Uii  ( .x(\U11/ni ), .a(i[11]) );
    inv_1 \U11/Uih  ( .x(\U11/nh ), .a(h[11]) );
    inv_1 \U11/Uil  ( .x(\U11/nl ), .a(l[11]) );
    ao23_1 \U11/Ucl/U1/U1  ( .x(l[11]), .a(n5), .b(l[11]), .c(n4), .d(\U11/ni 
        ), .e(\U11/nh ) );
    ao23_1 \U11/Uch/U1/U1  ( .x(h[11]), .a(n5), .b(h[11]), .c(n4), .d(i[11]), 
        .e(\U11/nl ) );
    inv_1 \U10/Uii  ( .x(\U10/ni ), .a(i[10]) );
    inv_1 \U10/Uih  ( .x(\U10/nh ), .a(h[10]) );
    inv_1 \U10/Uil  ( .x(\U10/nl ), .a(l[10]) );
    ao23_1 \U10/Ucl/U1/U1  ( .x(l[10]), .a(n5), .b(l[10]), .c(n3), .d(\U10/ni 
        ), .e(\U10/nh ) );
    ao23_1 \U10/Uch/U1/U1  ( .x(h[10]), .a(n5), .b(h[10]), .c(n3), .d(i[10]), 
        .e(\U10/nl ) );
    inv_1 \U9/Uii  ( .x(\U9/ni ), .a(i[9]) );
    inv_1 \U9/Uih  ( .x(\U9/nh ), .a(h[9]) );
    inv_1 \U9/Uil  ( .x(\U9/nl ), .a(l[9]) );
    ao23_1 \U9/Ucl/U1/U1  ( .x(l[9]), .a(n5), .b(l[9]), .c(n3), .d(\U9/ni ), 
        .e(\U9/nh ) );
    ao23_1 \U9/Uch/U1/U1  ( .x(h[9]), .a(n5), .b(h[9]), .c(n3), .d(i[9]), .e(
        \U9/nl ) );
    inv_1 \U8/Uii  ( .x(\U8/ni ), .a(i[8]) );
    inv_1 \U8/Uih  ( .x(\U8/nh ), .a(h[8]) );
    inv_1 \U8/Uil  ( .x(\U8/nl ), .a(l[8]) );
    ao23_1 \U8/Ucl/U1/U1  ( .x(l[8]), .a(n5), .b(l[8]), .c(n3), .d(\U8/ni ), 
        .e(\U8/nh ) );
    ao23_1 \U8/Uch/U1/U1  ( .x(h[8]), .a(n5), .b(h[8]), .c(n3), .d(i[8]), .e(
        \U8/nl ) );
    inv_1 \U7/Uii  ( .x(\U7/ni ), .a(i[7]) );
    inv_1 \U7/Uih  ( .x(\U7/nh ), .a(h[7]) );
    inv_1 \U7/Uil  ( .x(\U7/nl ), .a(l[7]) );
    ao23_1 \U7/Ucl/U1/U1  ( .x(l[7]), .a(n7), .b(l[7]), .c(n3), .d(\U7/ni ), 
        .e(\U7/nh ) );
    ao23_1 \U7/Uch/U1/U1  ( .x(h[7]), .a(n7), .b(h[7]), .c(n2), .d(i[7]), .e(
        \U7/nl ) );
    inv_1 \U6/Uii  ( .x(\U6/ni ), .a(i[6]) );
    inv_1 \U6/Uih  ( .x(\U6/nh ), .a(h[6]) );
    inv_1 \U6/Uil  ( .x(\U6/nl ), .a(l[6]) );
    ao23_1 \U6/Ucl/U1/U1  ( .x(l[6]), .a(n7), .b(l[6]), .c(n2), .d(\U6/ni ), 
        .e(\U6/nh ) );
    ao23_1 \U6/Uch/U1/U1  ( .x(h[6]), .a(n7), .b(h[6]), .c(n2), .d(i[6]), .e(
        \U6/nl ) );
    inv_1 \U5/Uii  ( .x(\U5/ni ), .a(i[5]) );
    inv_1 \U5/Uih  ( .x(\U5/nh ), .a(h[5]) );
    inv_1 \U5/Uil  ( .x(\U5/nl ), .a(l[5]) );
    ao23_1 \U5/Ucl/U1/U1  ( .x(l[5]), .a(n7), .b(l[5]), .c(n2), .d(\U5/ni ), 
        .e(\U5/nh ) );
    ao23_1 \U5/Uch/U1/U1  ( .x(h[5]), .a(n7), .b(h[5]), .c(n2), .d(i[5]), .e(
        \U5/nl ) );
    inv_1 \U4/Uii  ( .x(\U4/ni ), .a(i[4]) );
    inv_1 \U4/Uih  ( .x(\U4/nh ), .a(h[4]) );
    inv_1 \U4/Uil  ( .x(\U4/nl ), .a(l[4]) );
    ao23_1 \U4/Ucl/U1/U1  ( .x(l[4]), .a(n6), .b(l[4]), .c(n2), .d(\U4/ni ), 
        .e(\U4/nh ) );
    ao23_1 \U4/Uch/U1/U1  ( .x(h[4]), .a(n6), .b(h[4]), .c(n2), .d(i[4]), .e(
        \U4/nl ) );
    inv_1 \U3/Uii  ( .x(\U3/ni ), .a(i[3]) );
    inv_1 \U3/Uih  ( .x(\U3/nh ), .a(h[3]) );
    inv_1 \U3/Uil  ( .x(\U3/nl ), .a(l[3]) );
    ao23_1 \U3/Ucl/U1/U1  ( .x(l[3]), .a(n6), .b(l[3]), .c(n2), .d(\U3/ni ), 
        .e(\U3/nh ) );
    ao23_1 \U3/Uch/U1/U1  ( .x(h[3]), .a(n8), .b(h[3]), .c(n1), .d(i[3]), .e(
        \U3/nl ) );
    inv_1 \U2/Uii  ( .x(\U2/ni ), .a(i[2]) );
    inv_1 \U2/Uih  ( .x(\U2/nh ), .a(h[2]) );
    inv_1 \U2/Uil  ( .x(\U2/nl ), .a(l[2]) );
    ao23_1 \U2/Ucl/U1/U1  ( .x(l[2]), .a(n8), .b(l[2]), .c(n1), .d(\U2/ni ), 
        .e(\U2/nh ) );
    ao23_1 \U2/Uch/U1/U1  ( .x(h[2]), .a(n8), .b(h[2]), .c(n1), .d(i[2]), .e(
        \U2/nl ) );
    inv_1 \U1/Uii  ( .x(\U1/ni ), .a(i[1]) );
    inv_1 \U1/Uih  ( .x(\U1/nh ), .a(h[1]) );
    inv_1 \U1/Uil  ( .x(\U1/nl ), .a(l[1]) );
    ao23_1 \U1/Ucl/U1/U1  ( .x(l[1]), .a(n8), .b(l[1]), .c(n1), .d(\U1/ni ), 
        .e(\U1/nh ) );
    ao23_1 \U1/Uch/U1/U1  ( .x(h[1]), .a(n8), .b(h[1]), .c(n1), .d(i[1]), .e(
        \U1/nl ) );
    inv_1 \U0/Uii  ( .x(\U0/ni ), .a(i[0]) );
    inv_1 \U0/Uih  ( .x(\U0/nh ), .a(h[0]) );
    inv_1 \U0/Uil  ( .x(\U0/nl ), .a(l[0]) );
    ao23_1 \U0/Ucl/U1/U1  ( .x(l[0]), .a(n8), .b(l[0]), .c(n1), .d(\U0/ni ), 
        .e(\U0/nh ) );
    ao23_1 \U0/Uch/U1/U1  ( .x(h[0]), .a(n8), .b(h[0]), .c(n1), .d(i[0]), .e(
        \U0/nl ) );
    buf_16 U1 ( .x(n1), .a(n12) );
    buf_16 U2 ( .x(n2), .a(n12) );
    buf_16 U3 ( .x(n3), .a(n12) );
    buf_16 U4 ( .x(n4), .a(n11) );
    buf_16 U5 ( .x(n5), .a(n11) );
    buf_16 U6 ( .x(n6), .a(n11) );
    buf_16 U7 ( .x(n7), .a(n10) );
    buf_16 U8 ( .x(n8), .a(n10) );
    buf_16 U9 ( .x(n9), .a(n10) );
    buf_16 U10 ( .x(n10), .a(req) );
    buf_16 U11 ( .x(n11), .a(req) );
    buf_16 U12 ( .x(n12), .a(req) );
endmodule


module latch_ctrl_0 ( rin, ain, rout, aout, en, reset );
input  rin, aout, reset;
output ain, rout, en;
    wire N5, N6, na, a, n_rout, nreset, n3, \c_rout/ob , n1;
    inv_1 U0 ( .x(nreset), .a(reset) );
    nor2_1 U1 ( .x(ain), .a(na), .b(n1) );
    inv_1 U2 ( .x(na), .a(a) );
    inv_1 U3 ( .x(N6), .a(N5) );
    inv_1 U4 ( .x(rout), .a(n_rout) );
    and2_1 C9 ( .x(n3), .a(na), .b(N6) );
    or2_1 C11 ( .x(N5), .a(rout), .b(aout) );
    oa21_1 \c_na/__tmp99/U1  ( .x(a), .a(n1), .b(a), .c(rin) );
    oai21_1 \c_rout/U1  ( .x(\c_rout/ob ), .a(aout), .b(n_rout), .c(na) );
    nand2_1 \c_rout/U2  ( .x(n_rout), .a(nreset), .b(\c_rout/ob ) );
    buf_1 U5 ( .x(en), .a(n3) );
    buf_1 U6 ( .x(n1), .a(n3) );
endmodule


module m2cp_iport ( req_in, ts_o, sel_o, mult_o, we_o, prd_o, seq_o, adr_o, 
    dat_o, ain, ic_seq, ic_pred, ic_size, ic_itag, ic_wd, ic_lock, ic_a, 
    ic_rnw, ic_col, ic_ack, req_out, ts_i, we_i, err_i, rty_i, acc_i, dat_i, 
    aout, ir_rd, ir_err, ir_rnw, ir_ack, tag_id, reset );
input  [2:0] ts_o;
input  [3:0] sel_o;
input  [31:0] adr_o;
input  [31:0] dat_o;
output [1:0] ic_seq;
output [1:0] ic_pred;
output [3:0] ic_size;
output [9:0] ic_itag;
output [63:0] ic_wd;
output [1:0] ic_lock;
output [63:0] ic_a;
output [1:0] ic_rnw;
output [5:0] ic_col;
output [2:0] ts_i;
output [31:0] dat_i;
input  [63:0] ir_rd;
input  [1:0] ir_err;
input  [1:0] ir_rnw;
input  [4:0] tag_id;
input  req_in, mult_o, we_o, prd_o, seq_o, ic_ack, aout, reset;
output ain, req_out, we_i, err_i, rty_i, acc_i, ir_ack;
    wire n63, n64, n65, n68, n69, n70, n72, n73, n74, n75, n76, n77, n78, n79, 
        n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, 
        n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, 
        n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
        n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, 
        n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
        n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
        n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
        n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
        n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
        n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, 
        n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, 
        n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, 
        n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, 
        n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, 
        n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, 
        n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, 
        n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, 
        n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, 
        n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n2, n3, n4, 
        n5, req_in_delayed, \size[1] , \size[0] , \data[15] , \data[14] , 
        \data[13] , \data[12] , \data[11] , \data[10] , \data[9] , \data[8] , 
        \data[7] , \data[6] , \data[5] , \data[4] , \data[3] , \data[2] , 
        \data[1] , \data[0] , _24_net_, _25_net_, _26_net_, comp_basic, 
        high_ir_rd, low_ir_rd, comp_rd, _27_net_, all_r, _28_net_, all_w, 
        complete, complete_delayed, en, \all_read/__tmp99/loop , \Ucol2/nl , 
        \Ucol2/ni , \Ucol2/nh , \Ucol1/nl , \Ucol1/ni , \Ucol1/nh , \Ucol0/nl , 
        \Ucol0/ni , \Ucol0/nh , \Utag4/nl , \Utag4/ni , \Utag4/nh , \Utag3/nl , 
        \Utag3/ni , \Utag3/nh , \Utag2/nl , \Utag2/ni , \Utag2/nh , \Utag1/nl , 
        \Utag1/ni , \Utag1/nh , \Utag0/nl , \Utag0/ni , \Utag0/nh , \Usze1/nl , 
        \Usze1/ni , \Usze1/nh , \Usze0/nl , \Usze0/ni , \Usze0/nh , \Urnw/nl , 
        \Urnw/ni , \Urnw/nh , \Ulock/nl , \Ulock/ni , \Ulock/nh , \Upred/nl , 
        \Upred/ni , \Upred/nh , \Useq/nl , \Useq/ni , \Useq/nh , n1, n6, n7, 
        n8, n9, n10, n11;
    assign ain = ic_ack;
    assign ts_i[2] = 1'b0;
    assign ts_i[1] = 1'b0;
    assign ts_i[0] = 1'b0;
    assign rty_i = 1'b0;
    assign acc_i = 1'b0;
    matched_delay_m2cp_com_iport U130 ( .x(req_in_delayed), .a(req_in) );
    sr2dr_word_1 Uwd ( .i({dat_o[31], dat_o[30], dat_o[29], dat_o[28], 
        dat_o[27], dat_o[26], dat_o[25], dat_o[24], dat_o[23], dat_o[22], 
        dat_o[21], dat_o[20], dat_o[19], dat_o[18], dat_o[17], dat_o[16], 
        \data[15] , \data[14] , \data[13] , \data[12] , \data[11] , \data[10] , 
        \data[9] , \data[8] , \data[7] , \data[6] , \data[5] , \data[4] , 
        \data[3] , \data[2] , \data[1] , \data[0] }), .req(n8), .h(ic_wd
        [63:32]), .l(ic_wd[31:0]) );
    sr2dr_word_0 Ua ( .i(adr_o), .req(n8), .h(ic_a[63:32]), .l(ic_a[31:0]) );
    latch_ctrl_0 lc ( .rin(complete_delayed), .ain(ir_ack), .rout(req_out), 
        .aout(aout), .en(en), .reset(reset) );
    nand2_1 U61 ( .x(_26_net_), .a(n72), .b(n77) );
    and2_1 U274 ( .x(_27_net_), .a(ir_rnw[1]), .b(ir_err[0]) );
    inv_1 U275 ( .x(_24_net_), .a(we_o) );
    inv_1 U2 ( .x(n112), .a(ir_rd[4]) );
    inv_1 U3 ( .x(n124), .a(ir_rd[0]) );
    inv_1 U4 ( .x(n118), .a(ir_rd[2]) );
    inv_1 U5 ( .x(n206), .a(dat_o[28]) );
    inv_1 U6 ( .x(n208), .a(dat_o[27]) );
    inv_1 U7 ( .x(n210), .a(dat_o[26]) );
    inv_1 U8 ( .x(n197), .a(dat_o[25]) );
    inv_1 U9 ( .x(n199), .a(dat_o[24]) );
    inv_1 U10 ( .x(n202), .a(dat_o[15]) );
    inv_1 U11 ( .x(n201), .a(dat_o[31]) );
    inv_1 U12 ( .x(n203), .a(dat_o[30]) );
    inv_1 U13 ( .x(n204), .a(dat_o[29]) );
    nor2_1 U14 ( .x(\size[1] ), .a(n83), .b(n84) );
    inv_1 U15 ( .x(n72), .a(ir_rnw[0]) );
    oa21_1 U16 ( .x(n89), .a(n205), .b(n64), .c(n2) );
    inv_1 U24 ( .x(n2), .a(n90) );
    inv_1 U17 ( .x(n205), .a(dat_o[13]) );
    inv_1 U18 ( .x(n64), .a(sel_o[1]) );
    oa21_1 U19 ( .x(n97), .a(n198), .b(n64), .c(n3) );
    inv_1 U276 ( .x(n3), .a(n98) );
    inv_1 U20 ( .x(n198), .a(dat_o[9]) );
    oa21_1 U21 ( .x(n87), .a(n63), .b(n64), .c(n4) );
    inv_1 U277 ( .x(n4), .a(n88) );
    inv_1 U22 ( .x(n63), .a(dat_o[14]) );
    oa21_1 U23 ( .x(n85), .a(n202), .b(n64), .c(n5) );
    inv_1 U278 ( .x(n5), .a(n86) );
    nand2_1 U25 ( .x(n290), .a(n289), .b(n288) );
    nand2_1 U26 ( .x(n79), .a(n277), .b(n270) );
    nor2_1 U27 ( .x(n277), .a(n273), .b(n276) );
    nor2_1 U28 ( .x(n270), .a(n266), .b(n269) );
    nand2_1 U29 ( .x(n283), .a(n282), .b(n281) );
    nand2_1 U30 ( .x(n298), .a(dat_o[20]), .b(n70) );
    inv_1 U31 ( .x(n70), .a(n68) );
    nand2_1 U32 ( .x(n213), .a(n223), .b(sel_o[1]) );
    nand2_1 U33 ( .x(n80), .a(n291), .b(n284) );
    nor2_1 U34 ( .x(n291), .a(n287), .b(n290) );
    nor2_1 U35 ( .x(n284), .a(n280), .b(n283) );
    aoi21_1 U36 ( .x(n99), .a(dat_o[8]), .b(sel_o[1]), .c(n100) );
    aoi21_1 U37 ( .x(n95), .a(dat_o[10]), .b(sel_o[1]), .c(n96) );
    aoi21_1 U38 ( .x(n93), .a(dat_o[11]), .b(sel_o[1]), .c(n94) );
    aoi21_1 U39 ( .x(n91), .a(dat_o[12]), .b(sel_o[1]), .c(n92) );
    inv_1 U40 ( .x(n81), .a(all_r) );
    nand2_1 U42 ( .x(n84), .a(sel_o[0]), .b(sel_o[1]) );
    inv_1 U45 ( .x(n68), .a(sel_o[2]) );
    inv_1 U46 ( .x(n69), .a(n68) );
    nand2_1 U51 ( .x(n300), .a(dat_o[19]), .b(n69) );
    nand2_1 U52 ( .x(n294), .a(dat_o[22]), .b(n69) );
    nand2_1 U53 ( .x(n302), .a(dat_o[18]), .b(n69) );
    nand2_1 U54 ( .x(n296), .a(dat_o[21]), .b(n69) );
    nand2_1 U55 ( .x(n306), .a(dat_o[16]), .b(n69) );
    nand2_1 U56 ( .x(n292), .a(dat_o[23]), .b(n69) );
    nand2_1 U57 ( .x(n304), .a(dat_o[17]), .b(n69) );
    nand4_1 U60 ( .x(low_ir_rd), .a(n73), .b(n74), .c(n75), .d(n76) );
    nand2_1 U62 ( .x(complete), .a(n81), .b(n82) );
    matched_delay_m2cp_resp_iport mdel ( .x(complete_delayed), .a(complete) );
    inv_1 U63 ( .x(n200), .a(dat_o[8]) );
    inv_1 U64 ( .x(n207), .a(dat_o[12]) );
    inv_1 U65 ( .x(n209), .a(dat_o[11]) );
    inv_1 U66 ( .x(n211), .a(dat_o[10]) );
    nand4_1 U67 ( .x(n224), .a(n225), .b(n226), .c(n227), .d(n228) );
    nand4_1 U68 ( .x(n229), .a(n230), .b(n231), .c(n232), .d(n233) );
    nor2_1 U69 ( .x(n76), .a(n224), .b(n229) );
    nand4_1 U70 ( .x(n234), .a(n235), .b(n236), .c(n237), .d(n238) );
    nand4_1 U71 ( .x(n239), .a(n240), .b(n241), .c(n242), .d(n243) );
    nor2_1 U72 ( .x(n75), .a(n234), .b(n239) );
    nand4_1 U73 ( .x(n244), .a(n245), .b(n246), .c(n247), .d(n248) );
    nand4_1 U74 ( .x(n249), .a(n250), .b(n251), .c(n252), .d(n253) );
    nor2_1 U75 ( .x(n74), .a(n244), .b(n249) );
    nand4_1 U76 ( .x(n254), .a(n255), .b(n256), .c(n257), .d(n258) );
    nand4_1 U77 ( .x(n259), .a(n260), .b(n261), .c(n262), .d(n263) );
    nor2_1 U78 ( .x(n73), .a(n254), .b(n259) );
    nand2_1 U79 ( .x(n266), .a(n265), .b(n264) );
    nand2_1 U80 ( .x(n269), .a(n268), .b(n267) );
    nand2_1 U81 ( .x(n273), .a(n272), .b(n271) );
    nand2_1 U82 ( .x(n276), .a(n275), .b(n274) );
    nand2_1 U83 ( .x(n280), .a(n279), .b(n278) );
    nand2_1 U84 ( .x(n287), .a(n286), .b(n285) );
    nand2_1 U85 ( .x(n86), .a(n292), .b(n293) );
    nand2_1 U86 ( .x(n88), .a(n294), .b(n295) );
    nand2_1 U87 ( .x(n90), .a(n296), .b(n297) );
    nand2_1 U88 ( .x(n92), .a(n298), .b(n299) );
    nand2_1 U89 ( .x(n94), .a(n300), .b(n301) );
    nand2_1 U90 ( .x(n96), .a(n302), .b(n303) );
    nand2_1 U91 ( .x(n98), .a(n304), .b(n305) );
    nand2_1 U92 ( .x(n100), .a(n306), .b(n307) );
    inv_1 U93 ( .x(n222), .a(dat_o[0]) );
    inv_1 U94 ( .x(n221), .a(dat_o[1]) );
    inv_1 U95 ( .x(n220), .a(dat_o[2]) );
    inv_1 U96 ( .x(n219), .a(dat_o[3]) );
    inv_1 U97 ( .x(n218), .a(dat_o[4]) );
    inv_1 U98 ( .x(n217), .a(dat_o[5]) );
    inv_1 U99 ( .x(n216), .a(dat_o[6]) );
    inv_1 U100 ( .x(n215), .a(dat_o[7]) );
    inv_1 U101 ( .x(n77), .a(ir_rnw[1]) );
    inv_1 U103 ( .x(n82), .a(all_w) );
    nand2_1 U104 ( .x(n293), .a(dat_o[31]), .b(sel_o[3]) );
    nand2_1 U105 ( .x(n295), .a(dat_o[30]), .b(sel_o[3]) );
    nand2_1 U109 ( .x(n303), .a(dat_o[26]), .b(sel_o[3]) );
    nand2_1 U110 ( .x(n305), .a(dat_o[25]), .b(sel_o[3]) );
    nand2_1 U111 ( .x(n307), .a(dat_o[24]), .b(sel_o[3]) );
    mux2i_1 U113 ( .x(\data[0] ), .d0(n99), .sl(n65), .d1(n222) );
    mux2i_1 U114 ( .x(\data[10] ), .d0(n211), .sl(n214), .d1(n210) );
    mux2i_1 U115 ( .x(\data[11] ), .d0(n209), .sl(n214), .d1(n208) );
    mux2i_1 U116 ( .x(\data[12] ), .d0(n207), .sl(n214), .d1(n206) );
    mux2i_1 U117 ( .x(\data[13] ), .d0(n205), .sl(n214), .d1(n204) );
    mux2i_1 U118 ( .x(\data[14] ), .d0(n63), .sl(n214), .d1(n203) );
    mux2i_1 U119 ( .x(\data[15] ), .d0(n202), .sl(n214), .d1(n201) );
    mux2i_1 U120 ( .x(\data[1] ), .d0(n97), .sl(n65), .d1(n221) );
    mux2i_1 U121 ( .x(\data[2] ), .d0(n95), .sl(n65), .d1(n220) );
    mux2i_1 U122 ( .x(\data[3] ), .d0(n93), .sl(n65), .d1(n219) );
    mux2i_1 U123 ( .x(\data[4] ), .d0(n91), .sl(n65), .d1(n218) );
    mux2i_1 U124 ( .x(\data[5] ), .d0(n89), .sl(n65), .d1(n217) );
    mux2i_1 U125 ( .x(\data[6] ), .d0(n87), .sl(n65), .d1(n216) );
    mux2i_1 U126 ( .x(\data[7] ), .d0(n85), .sl(n65), .d1(n215) );
    mux2i_1 U127 ( .x(\data[8] ), .d0(n200), .sl(n214), .d1(n199) );
    mux2i_1 U128 ( .x(\data[9] ), .d0(n198), .sl(n214), .d1(n197) );
    nor2_1 U129 ( .x(high_ir_rd), .a(n79), .b(n80) );
    mux2i_1 U131 ( .x(\size[0] ), .d0(n212), .sl(n65), .d1(n213) );
    nand2i_1 U132 ( .x(n308), .a(sel_o[1]), .b(n70) );
    inv_1 U133 ( .x(n255), .a(n182) );
    inv_1 U134 ( .x(n256), .a(n179) );
    inv_1 U135 ( .x(n257), .a(n176) );
    inv_1 U136 ( .x(n258), .a(n173) );
    inv_1 U137 ( .x(n260), .a(n194) );
    inv_1 U138 ( .x(n261), .a(n191) );
    inv_1 U139 ( .x(n262), .a(n188) );
    inv_1 U140 ( .x(n263), .a(n185) );
    inv_1 U141 ( .x(n245), .a(n158) );
    inv_1 U142 ( .x(n246), .a(n155) );
    inv_1 U143 ( .x(n247), .a(n152) );
    inv_1 U144 ( .x(n248), .a(n149) );
    inv_1 U145 ( .x(n250), .a(n170) );
    inv_1 U146 ( .x(n251), .a(n167) );
    inv_1 U147 ( .x(n252), .a(n164) );
    inv_1 U148 ( .x(n253), .a(n161) );
    inv_1 U149 ( .x(n235), .a(n134) );
    inv_1 U150 ( .x(n236), .a(n131) );
    inv_1 U151 ( .x(n237), .a(n128) );
    inv_1 U152 ( .x(n238), .a(n125) );
    inv_1 U153 ( .x(n240), .a(n146) );
    inv_1 U154 ( .x(n241), .a(n143) );
    inv_1 U155 ( .x(n242), .a(n140) );
    inv_1 U156 ( .x(n243), .a(n137) );
    inv_1 U157 ( .x(n225), .a(n110) );
    inv_1 U158 ( .x(n226), .a(n107) );
    inv_1 U159 ( .x(n227), .a(n104) );
    inv_1 U160 ( .x(n228), .a(n101) );
    inv_1 U161 ( .x(n230), .a(n122) );
    inv_1 U162 ( .x(n231), .a(n119) );
    inv_1 U163 ( .x(n232), .a(n116) );
    inv_1 U164 ( .x(n233), .a(n113) );
    nor2_1 U165 ( .x(n272), .a(n252), .b(n253) );
    nor2_1 U166 ( .x(n271), .a(n250), .b(n251) );
    nor2_1 U167 ( .x(n275), .a(n247), .b(n248) );
    nor2_1 U168 ( .x(n274), .a(n245), .b(n246) );
    nor2_1 U169 ( .x(n265), .a(n262), .b(n263) );
    nor2_1 U170 ( .x(n264), .a(n260), .b(n261) );
    nor2_1 U171 ( .x(n268), .a(n257), .b(n258) );
    nor2_1 U172 ( .x(n267), .a(n255), .b(n256) );
    nor2_1 U173 ( .x(n286), .a(n232), .b(n233) );
    nor2_1 U174 ( .x(n285), .a(n230), .b(n231) );
    nor2_1 U175 ( .x(n289), .a(n227), .b(n228) );
    nor2_1 U176 ( .x(n288), .a(n225), .b(n226) );
    nor2_1 U177 ( .x(n279), .a(n242), .b(n243) );
    nor2_1 U178 ( .x(n278), .a(n240), .b(n241) );
    nor2_1 U179 ( .x(n282), .a(n237), .b(n238) );
    nor2_1 U180 ( .x(n281), .a(n235), .b(n236) );
    nand2_1 U181 ( .x(n182), .a(n183), .b(n184) );
    nand2_1 U182 ( .x(n179), .a(n180), .b(n181) );
    nand2_1 U183 ( .x(n176), .a(n177), .b(n178) );
    nand2_1 U184 ( .x(n173), .a(n174), .b(n175) );
    nand2_1 U185 ( .x(n194), .a(n195), .b(n196) );
    nand2_1 U186 ( .x(n191), .a(n192), .b(n193) );
    nand2_1 U187 ( .x(n188), .a(n189), .b(n190) );
    nand2_1 U188 ( .x(n185), .a(n186), .b(n187) );
    nand2_1 U189 ( .x(n158), .a(n159), .b(n160) );
    nand2_1 U190 ( .x(n155), .a(n156), .b(n157) );
    nand2_1 U191 ( .x(n152), .a(n153), .b(n154) );
    nand2_1 U192 ( .x(n149), .a(n150), .b(n151) );
    nand2_1 U193 ( .x(n170), .a(n171), .b(n172) );
    nand2_1 U194 ( .x(n167), .a(n168), .b(n169) );
    nand2_1 U195 ( .x(n164), .a(n165), .b(n166) );
    nand2_1 U196 ( .x(n161), .a(n162), .b(n163) );
    nand2_1 U197 ( .x(n134), .a(n135), .b(n136) );
    nand2_1 U198 ( .x(n131), .a(n132), .b(n133) );
    nand2_1 U199 ( .x(n128), .a(n129), .b(n130) );
    nand2_1 U200 ( .x(n125), .a(n126), .b(n127) );
    nand2_1 U201 ( .x(n146), .a(n147), .b(n148) );
    nand2_1 U202 ( .x(n143), .a(n144), .b(n145) );
    nand2_1 U203 ( .x(n140), .a(n141), .b(n142) );
    nand2_1 U204 ( .x(n137), .a(n138), .b(n139) );
    nand2_1 U205 ( .x(n110), .a(n111), .b(n112) );
    nand2_1 U206 ( .x(n107), .a(n108), .b(n109) );
    nand2_1 U207 ( .x(n104), .a(n105), .b(n106) );
    nand2_1 U208 ( .x(n101), .a(n102), .b(n103) );
    nand2_1 U209 ( .x(n122), .a(n123), .b(n124) );
    nand2_1 U210 ( .x(n119), .a(n120), .b(n121) );
    nand2_1 U211 ( .x(n116), .a(n117), .b(n118) );
    nand2_1 U212 ( .x(n113), .a(n114), .b(n115) );
    inv_1 U213 ( .x(n183), .a(ir_rd[60]) );
    inv_1 U214 ( .x(n184), .a(ir_rd[28]) );
    inv_1 U215 ( .x(n180), .a(ir_rd[61]) );
    inv_1 U216 ( .x(n181), .a(ir_rd[29]) );
    inv_1 U217 ( .x(n177), .a(ir_rd[62]) );
    inv_1 U218 ( .x(n178), .a(ir_rd[30]) );
    inv_1 U219 ( .x(n174), .a(ir_rd[63]) );
    inv_1 U220 ( .x(n175), .a(ir_rd[31]) );
    inv_1 U221 ( .x(n195), .a(ir_rd[56]) );
    inv_1 U222 ( .x(n196), .a(ir_rd[24]) );
    inv_1 U223 ( .x(n192), .a(ir_rd[57]) );
    inv_1 U224 ( .x(n193), .a(ir_rd[25]) );
    inv_1 U225 ( .x(n189), .a(ir_rd[58]) );
    inv_1 U226 ( .x(n190), .a(ir_rd[26]) );
    inv_1 U227 ( .x(n186), .a(ir_rd[59]) );
    inv_1 U228 ( .x(n187), .a(ir_rd[27]) );
    inv_1 U229 ( .x(n159), .a(ir_rd[52]) );
    inv_1 U230 ( .x(n160), .a(ir_rd[20]) );
    inv_1 U231 ( .x(n156), .a(ir_rd[53]) );
    inv_1 U232 ( .x(n157), .a(ir_rd[21]) );
    inv_1 U233 ( .x(n153), .a(ir_rd[54]) );
    inv_1 U234 ( .x(n154), .a(ir_rd[22]) );
    inv_1 U235 ( .x(n150), .a(ir_rd[55]) );
    inv_1 U236 ( .x(n151), .a(ir_rd[23]) );
    inv_1 U237 ( .x(n171), .a(ir_rd[48]) );
    inv_1 U238 ( .x(n172), .a(ir_rd[16]) );
    inv_1 U239 ( .x(n168), .a(ir_rd[49]) );
    inv_1 U240 ( .x(n169), .a(ir_rd[17]) );
    inv_1 U241 ( .x(n165), .a(ir_rd[50]) );
    inv_1 U242 ( .x(n166), .a(ir_rd[18]) );
    inv_1 U243 ( .x(n162), .a(ir_rd[51]) );
    inv_1 U244 ( .x(n163), .a(ir_rd[19]) );
    inv_1 U245 ( .x(n135), .a(ir_rd[44]) );
    inv_1 U246 ( .x(n136), .a(ir_rd[12]) );
    inv_1 U247 ( .x(n132), .a(ir_rd[45]) );
    inv_1 U248 ( .x(n133), .a(ir_rd[13]) );
    inv_1 U249 ( .x(n129), .a(ir_rd[46]) );
    inv_1 U250 ( .x(n130), .a(ir_rd[14]) );
    inv_1 U251 ( .x(n126), .a(ir_rd[47]) );
    inv_1 U252 ( .x(n127), .a(ir_rd[15]) );
    inv_1 U253 ( .x(n147), .a(ir_rd[40]) );
    inv_1 U254 ( .x(n148), .a(ir_rd[8]) );
    inv_1 U255 ( .x(n144), .a(ir_rd[41]) );
    inv_1 U256 ( .x(n145), .a(ir_rd[9]) );
    inv_1 U257 ( .x(n141), .a(ir_rd[42]) );
    inv_1 U258 ( .x(n142), .a(ir_rd[10]) );
    inv_1 U259 ( .x(n138), .a(ir_rd[43]) );
    inv_1 U260 ( .x(n139), .a(ir_rd[11]) );
    inv_1 U261 ( .x(n111), .a(ir_rd[36]) );
    inv_1 U262 ( .x(n108), .a(ir_rd[37]) );
    inv_1 U263 ( .x(n109), .a(ir_rd[5]) );
    inv_1 U264 ( .x(n105), .a(ir_rd[38]) );
    inv_1 U265 ( .x(n106), .a(ir_rd[6]) );
    inv_1 U266 ( .x(n102), .a(ir_rd[39]) );
    inv_1 U267 ( .x(n103), .a(ir_rd[7]) );
    inv_1 U268 ( .x(n123), .a(ir_rd[32]) );
    inv_1 U269 ( .x(n120), .a(ir_rd[33]) );
    inv_1 U270 ( .x(n121), .a(ir_rd[1]) );
    inv_1 U271 ( .x(n117), .a(ir_rd[34]) );
    inv_1 U272 ( .x(n114), .a(ir_rd[35]) );
    inv_1 U273 ( .x(n115), .a(ir_rd[3]) );
    latn_1 \dat_i_reg[30]  ( .q(dat_i[30]), .d(ir_rd[62]), .g(n7) );
    latn_1 \dat_i_reg[28]  ( .q(dat_i[28]), .d(ir_rd[60]), .g(n7) );
    latn_1 \dat_i_reg[27]  ( .q(dat_i[27]), .d(ir_rd[59]), .g(n7) );
    latn_1 \dat_i_reg[26]  ( .q(dat_i[26]), .d(ir_rd[58]), .g(n7) );
    latn_1 \dat_i_reg[25]  ( .q(dat_i[25]), .d(ir_rd[57]), .g(n7) );
    latn_1 \dat_i_reg[24]  ( .q(dat_i[24]), .d(ir_rd[56]), .g(n7) );
    latn_1 \dat_i_reg[22]  ( .q(dat_i[22]), .d(ir_rd[54]), .g(n7) );
    latn_1 \dat_i_reg[20]  ( .q(dat_i[20]), .d(ir_rd[52]), .g(n7) );
    latn_1 \dat_i_reg[19]  ( .q(dat_i[19]), .d(ir_rd[51]), .g(n7) );
    latn_1 \dat_i_reg[18]  ( .q(dat_i[18]), .d(ir_rd[50]), .g(n7) );
    latn_1 \dat_i_reg[17]  ( .q(dat_i[17]), .d(ir_rd[49]), .g(n7) );
    latn_1 \dat_i_reg[16]  ( .q(dat_i[16]), .d(ir_rd[48]), .g(n6) );
    latn_1 \dat_i_reg[14]  ( .q(dat_i[14]), .d(ir_rd[46]), .g(n6) );
    latn_1 \dat_i_reg[12]  ( .q(dat_i[12]), .d(ir_rd[44]), .g(n6) );
    latn_1 \dat_i_reg[10]  ( .q(dat_i[10]), .d(ir_rd[42]), .g(n6) );
    latn_1 \dat_i_reg[8]  ( .q(dat_i[8]), .d(ir_rd[40]), .g(n6) );
    latn_1 \dat_i_reg[6]  ( .q(dat_i[6]), .d(ir_rd[38]), .g(n6) );
    latn_1 \dat_i_reg[4]  ( .q(dat_i[4]), .d(ir_rd[36]), .g(n6) );
    latn_1 \dat_i_reg[3]  ( .q(dat_i[3]), .d(ir_rd[35]), .g(n1) );
    latn_1 \dat_i_reg[2]  ( .q(dat_i[2]), .d(ir_rd[34]), .g(n1) );
    latn_1 \dat_i_reg[1]  ( .q(dat_i[1]), .d(ir_rd[33]), .g(n1) );
    latn_1 \dat_i_reg[0]  ( .q(dat_i[0]), .d(ir_rd[32]), .g(n1) );
    latn_1 we_i_reg ( .q(we_i), .d(ir_rnw[0]), .g(n1) );
    latn_1 err_i_reg ( .q(err_i), .d(ir_err[1]), .g(n1) );
    latn_1 \dat_i_reg[13]  ( .q(dat_i[13]), .d(ir_rd[45]), .g(n6) );
    latn_1 \dat_i_reg[5]  ( .q(dat_i[5]), .d(ir_rd[37]), .g(n1) );
    latn_1 \dat_i_reg[15]  ( .q(dat_i[15]), .d(ir_rd[47]), .g(n6) );
    latn_1 \dat_i_reg[7]  ( .q(dat_i[7]), .d(ir_rd[39]), .g(n1) );
    latn_1 \dat_i_reg[29]  ( .q(dat_i[29]), .d(ir_rd[61]), .g(n6) );
    latn_1 \dat_i_reg[21]  ( .q(dat_i[21]), .d(ir_rd[53]), .g(n1) );
    latn_1 \dat_i_reg[31]  ( .q(dat_i[31]), .d(ir_rd[63]), .g(n6) );
    latn_1 \dat_i_reg[23]  ( .q(dat_i[23]), .d(ir_rd[55]), .g(n1) );
    latn_1 \dat_i_reg[9]  ( .q(dat_i[9]), .d(ir_rd[41]), .g(n6) );
    latn_1 \dat_i_reg[11]  ( .q(dat_i[11]), .d(ir_rd[43]), .g(n1) );
    oa21_1 \all_write/__tmp99/U1  ( .x(all_w), .a(_28_net_), .b(all_w), .c(
        comp_basic) );
    ao31_1 \all_read/__tmp99/aoi  ( .x(\all_read/__tmp99/loop ), .a(comp_basic
        ), .b(comp_rd), .c(_27_net_), .d(all_r) );
    oa21_1 \all_read/__tmp99/outGate  ( .x(all_r), .a(comp_basic), .b(comp_rd), 
        .c(\all_read/__tmp99/loop ) );
    ao222_1 \rd/__tmp99/U1  ( .x(comp_rd), .a(high_ir_rd), .b(low_ir_rd), .c(
        high_ir_rd), .d(comp_rd), .e(low_ir_rd), .f(comp_rd) );
    ao222_1 \basic/__tmp99/U1  ( .x(comp_basic), .a(_25_net_), .b(_26_net_), 
        .c(_25_net_), .d(comp_basic), .e(_26_net_), .f(comp_basic) );
    inv_1 \Ucol2/Uii  ( .x(\Ucol2/ni ), .a(ts_o[2]) );
    inv_1 \Ucol2/Uih  ( .x(\Ucol2/nh ), .a(ic_col[5]) );
    inv_1 \Ucol2/Uil  ( .x(\Ucol2/nl ), .a(ic_col[2]) );
    ao23_1 \Ucol2/Ucl/U1/U1  ( .x(ic_col[2]), .a(n11), .b(ic_col[2]), .c(n8), 
        .d(\Ucol2/ni ), .e(\Ucol2/nh ) );
    ao23_1 \Ucol2/Uch/U1/U1  ( .x(ic_col[5]), .a(n11), .b(ic_col[5]), .c(n8), 
        .d(ts_o[2]), .e(\Ucol2/nl ) );
    inv_1 \Ucol1/Uii  ( .x(\Ucol1/ni ), .a(ts_o[1]) );
    inv_1 \Ucol1/Uih  ( .x(\Ucol1/nh ), .a(ic_col[4]) );
    inv_1 \Ucol1/Uil  ( .x(\Ucol1/nl ), .a(ic_col[1]) );
    ao23_1 \Ucol1/Ucl/U1/U1  ( .x(ic_col[1]), .a(n11), .b(ic_col[1]), .c(n8), 
        .d(\Ucol1/ni ), .e(\Ucol1/nh ) );
    ao23_1 \Ucol1/Uch/U1/U1  ( .x(ic_col[4]), .a(n11), .b(ic_col[4]), .c(n9), 
        .d(ts_o[1]), .e(\Ucol1/nl ) );
    inv_1 \Ucol0/Uii  ( .x(\Ucol0/ni ), .a(ts_o[0]) );
    inv_1 \Ucol0/Uih  ( .x(\Ucol0/nh ), .a(ic_col[3]) );
    inv_1 \Ucol0/Uil  ( .x(\Ucol0/nl ), .a(ic_col[0]) );
    ao23_1 \Ucol0/Ucl/U1/U1  ( .x(ic_col[0]), .a(n11), .b(ic_col[0]), .c(n10), 
        .d(\Ucol0/ni ), .e(\Ucol0/nh ) );
    ao23_1 \Ucol0/Uch/U1/U1  ( .x(ic_col[3]), .a(n11), .b(ic_col[3]), .c(n9), 
        .d(ts_o[0]), .e(\Ucol0/nl ) );
    inv_1 \Utag4/Uii  ( .x(\Utag4/ni ), .a(tag_id[4]) );
    inv_1 \Utag4/Uih  ( .x(\Utag4/nh ), .a(ic_itag[9]) );
    inv_1 \Utag4/Uil  ( .x(\Utag4/nl ), .a(ic_itag[4]) );
    ao23_1 \Utag4/Ucl/U1/U1  ( .x(ic_itag[4]), .a(n11), .b(ic_itag[4]), .c(n9), 
        .d(\Utag4/ni ), .e(\Utag4/nh ) );
    ao23_1 \Utag4/Uch/U1/U1  ( .x(ic_itag[9]), .a(n10), .b(ic_itag[9]), .c(n9), 
        .d(tag_id[4]), .e(\Utag4/nl ) );
    inv_1 \Utag3/Uii  ( .x(\Utag3/ni ), .a(tag_id[3]) );
    inv_1 \Utag3/Uih  ( .x(\Utag3/nh ), .a(ic_itag[8]) );
    inv_1 \Utag3/Uil  ( .x(\Utag3/nl ), .a(ic_itag[3]) );
    ao23_1 \Utag3/Ucl/U1/U1  ( .x(ic_itag[3]), .a(n10), .b(ic_itag[3]), .c(n9), 
        .d(\Utag3/ni ), .e(\Utag3/nh ) );
    ao23_1 \Utag3/Uch/U1/U1  ( .x(ic_itag[8]), .a(n10), .b(ic_itag[8]), .c(n9), 
        .d(tag_id[3]), .e(\Utag3/nl ) );
    inv_1 \Utag2/Uii  ( .x(\Utag2/ni ), .a(tag_id[2]) );
    inv_1 \Utag2/Uih  ( .x(\Utag2/nh ), .a(ic_itag[7]) );
    inv_1 \Utag2/Uil  ( .x(\Utag2/nl ), .a(ic_itag[2]) );
    ao23_1 \Utag2/Ucl/U1/U1  ( .x(ic_itag[2]), .a(n10), .b(ic_itag[2]), .c(n9), 
        .d(\Utag2/ni ), .e(\Utag2/nh ) );
    ao23_1 \Utag2/Uch/U1/U1  ( .x(ic_itag[7]), .a(n10), .b(ic_itag[7]), .c(n10
        ), .d(tag_id[2]), .e(\Utag2/nl ) );
    inv_1 \Utag1/Uii  ( .x(\Utag1/ni ), .a(tag_id[1]) );
    inv_1 \Utag1/Uih  ( .x(\Utag1/nh ), .a(ic_itag[6]) );
    inv_1 \Utag1/Uil  ( .x(\Utag1/nl ), .a(ic_itag[1]) );
    ao23_1 \Utag1/Ucl/U1/U1  ( .x(ic_itag[1]), .a(n11), .b(ic_itag[1]), .c(n9), 
        .d(\Utag1/ni ), .e(\Utag1/nh ) );
    ao23_1 \Utag1/Uch/U1/U1  ( .x(ic_itag[6]), .a(n11), .b(ic_itag[6]), .c(n9), 
        .d(tag_id[1]), .e(\Utag1/nl ) );
    inv_1 \Utag0/Uii  ( .x(\Utag0/ni ), .a(tag_id[0]) );
    inv_1 \Utag0/Uih  ( .x(\Utag0/nh ), .a(ic_itag[5]) );
    inv_1 \Utag0/Uil  ( .x(\Utag0/nl ), .a(ic_itag[0]) );
    ao23_1 \Utag0/Ucl/U1/U1  ( .x(ic_itag[0]), .a(n11), .b(ic_itag[0]), .c(n8), 
        .d(\Utag0/ni ), .e(\Utag0/nh ) );
    ao23_1 \Utag0/Uch/U1/U1  ( .x(ic_itag[5]), .a(n10), .b(ic_itag[5]), .c(n8), 
        .d(tag_id[0]), .e(\Utag0/nl ) );
    inv_1 \Usze1/Uii  ( .x(\Usze1/ni ), .a(\size[1] ) );
    inv_1 \Usze1/Uih  ( .x(\Usze1/nh ), .a(ic_size[3]) );
    inv_1 \Usze1/Uil  ( .x(\Usze1/nl ), .a(ic_size[1]) );
    ao23_1 \Usze1/Ucl/U1/U1  ( .x(ic_size[1]), .a(n10), .b(ic_size[1]), .c(n9), 
        .d(\Usze1/ni ), .e(\Usze1/nh ) );
    ao23_1 \Usze1/Uch/U1/U1  ( .x(ic_size[3]), .a(n10), .b(ic_size[3]), .c(n9), 
        .d(\size[1] ), .e(\Usze1/nl ) );
    inv_1 \Usze0/Uii  ( .x(\Usze0/ni ), .a(\size[0] ) );
    inv_1 \Usze0/Uih  ( .x(\Usze0/nh ), .a(ic_size[2]) );
    inv_1 \Usze0/Uil  ( .x(\Usze0/nl ), .a(ic_size[0]) );
    ao23_1 \Usze0/Ucl/U1/U1  ( .x(ic_size[0]), .a(n10), .b(ic_size[0]), .c(n9), 
        .d(\Usze0/ni ), .e(\Usze0/nh ) );
    ao23_1 \Usze0/Uch/U1/U1  ( .x(ic_size[2]), .a(n10), .b(ic_size[2]), .c(n9), 
        .d(\size[0] ), .e(\Usze0/nl ) );
    inv_1 \Urnw/Uii  ( .x(\Urnw/ni ), .a(_24_net_) );
    inv_1 \Urnw/Uih  ( .x(\Urnw/nh ), .a(ic_rnw[1]) );
    inv_1 \Urnw/Uil  ( .x(\Urnw/nl ), .a(ic_rnw[0]) );
    ao23_1 \Urnw/Ucl/U1/U1  ( .x(ic_rnw[0]), .a(n10), .b(ic_rnw[0]), .c(n9), 
        .d(\Urnw/ni ), .e(\Urnw/nh ) );
    ao23_1 \Urnw/Uch/U1/U1  ( .x(ic_rnw[1]), .a(n10), .b(ic_rnw[1]), .c(n9), 
        .d(_24_net_), .e(\Urnw/nl ) );
    inv_1 \Ulock/Uii  ( .x(\Ulock/ni ), .a(mult_o) );
    inv_1 \Ulock/Uih  ( .x(\Ulock/nh ), .a(ic_lock[1]) );
    inv_1 \Ulock/Uil  ( .x(\Ulock/nl ), .a(ic_lock[0]) );
    ao23_1 \Ulock/Ucl/U1/U1  ( .x(ic_lock[0]), .a(n11), .b(ic_lock[0]), .c(n9), 
        .d(\Ulock/ni ), .e(\Ulock/nh ) );
    ao23_1 \Ulock/Uch/U1/U1  ( .x(ic_lock[1]), .a(n11), .b(ic_lock[1]), .c(n8), 
        .d(mult_o), .e(\Ulock/nl ) );
    inv_1 \Upred/Uii  ( .x(\Upred/ni ), .a(prd_o) );
    inv_1 \Upred/Uih  ( .x(\Upred/nh ), .a(ic_pred[1]) );
    inv_1 \Upred/Uil  ( .x(\Upred/nl ), .a(ic_pred[0]) );
    ao23_1 \Upred/Ucl/U1/U1  ( .x(ic_pred[0]), .a(n11), .b(ic_pred[0]), .c(n8), 
        .d(\Upred/ni ), .e(\Upred/nh ) );
    ao23_1 \Upred/Uch/U1/U1  ( .x(ic_pred[1]), .a(n10), .b(ic_pred[1]), .c(n8), 
        .d(prd_o), .e(\Upred/nl ) );
    inv_1 \Useq/Uii  ( .x(\Useq/ni ), .a(seq_o) );
    inv_1 \Useq/Uih  ( .x(\Useq/nh ), .a(ic_seq[1]) );
    inv_1 \Useq/Uil  ( .x(\Useq/nl ), .a(ic_seq[0]) );
    ao23_1 \Useq/Ucl/U1/U1  ( .x(ic_seq[0]), .a(n10), .b(ic_seq[0]), .c(n8), 
        .d(\Useq/ni ), .e(\Useq/nh ) );
    ao23_1 \Useq/Uch/U1/U1  ( .x(ic_seq[1]), .a(n11), .b(ic_seq[1]), .c(n8), 
        .d(seq_o), .e(\Useq/nl ) );
    buf_3 U1 ( .x(n1), .a(en) );
    buf_3 U41 ( .x(n7), .a(en) );
    buf_3 U43 ( .x(n6), .a(en) );
    inv_2 U44 ( .x(n214), .a(n308) );
    buf_3 U47 ( .x(n65), .a(sel_o[0]) );
    nand3i_0 U48 ( .x(n212), .a(sel_o[1]), .b(sel_o[3]), .c(n70) );
    nor2_0 U49 ( .x(n223), .a(n70), .b(sel_o[3]) );
    nand2_0 U50 ( .x(n297), .a(dat_o[29]), .b(sel_o[3]) );
    nand2_0 U58 ( .x(n301), .a(dat_o[27]), .b(sel_o[3]) );
    nand2_0 U59 ( .x(n299), .a(dat_o[28]), .b(sel_o[3]) );
    nand2_0 U102 ( .x(n83), .a(n70), .b(sel_o[3]) );
    inv_0 U106 ( .x(n78), .a(ir_err[0]) );
    nand2i_0 U107 ( .x(_28_net_), .a(ir_err[1]), .b(n72) );
    nand2i_0 U108 ( .x(_25_net_), .a(ir_err[1]), .b(n78) );
    buf_16 U112 ( .x(n8), .a(req_in_delayed) );
    buf_16 U279 ( .x(n9), .a(req_in_delayed) );
    buf_16 U280 ( .x(n10), .a(req_in_delayed) );
    buf_16 U281 ( .x(n11), .a(req_in_delayed) );
endmodule


module master_if_iport ( nReset, mc_req, mc_we, mc_mult, mc_prd, mc_seq, mc_ts, 
    mc_sel, mc_adr, mc_dat, mc_ack, mr_req, mr_we, mr_err, mr_rty, mr_acc, 
    mr_ts, mr_sel, mr_dat, mr_ack, chaincommand, nchaincommandack, 
    chainresponse, nchainresponseack, e_bare, e_dm, e_im, e_wish, r_bare, r_dm, 
    r_im, r_wish, tag_id, force_bare );
input  [2:0] mc_ts;
input  [3:0] mc_sel;
input  [31:0] mc_adr;
input  [31:0] mc_dat;
output [2:0] mr_ts;
output [3:0] mr_sel;
output [31:0] mr_dat;
output [4:0] chaincommand;
input  [4:0] chainresponse;
input  [3:0] e_bare;
input  [3:0] e_dm;
input  [3:0] e_im;
input  [3:0] e_wish;
input  [3:0] r_bare;
input  [3:0] r_dm;
input  [3:0] r_im;
input  [3:0] r_wish;
input  [4:0] tag_id;
input  nReset, mc_req, mc_we, mc_mult, mc_prd, mc_seq, mr_ack, 
    nchaincommandack, force_bare;
output mc_ack, mr_req, mr_we, mr_err, mr_rty, mr_acc, nchainresponseack;
    wire \ci_seq[1] , \ci_seq[0] , \ci_lock[1] , \ci_lock[0] , \ci_rnw[1] , 
        \ci_rnw[0] , \ci_size[3] , \ci_size[2] , \ci_size[1] , \ci_size[0] , 
        \ci_itag[9] , \ci_itag[8] , \ci_itag[7] , \ci_itag[6] , \ci_itag[5] , 
        \ci_itag[4] , \ci_itag[3] , \ci_itag[2] , \ci_itag[1] , \ci_itag[0] , 
        \ci_a[63] , \ci_a[62] , \ci_a[61] , \ci_a[60] , \ci_a[59] , \ci_a[58] , 
        \ci_a[57] , \ci_a[56] , \ci_a[55] , \ci_a[54] , \ci_a[53] , \ci_a[52] , 
        \ci_a[51] , \ci_a[50] , \ci_a[49] , \ci_a[48] , \ci_a[47] , \ci_a[46] , 
        \ci_a[45] , \ci_a[44] , \ci_a[43] , \ci_a[42] , \ci_a[41] , \ci_a[40] , 
        \ci_a[39] , \ci_a[38] , \ci_a[37] , \ci_a[36] , \ci_a[35] , \ci_a[34] , 
        \ci_a[33] , \ci_a[32] , \ci_a[31] , \ci_a[30] , \ci_a[29] , \ci_a[28] , 
        \ci_a[27] , \ci_a[26] , \ci_a[25] , \ci_a[24] , \ci_a[23] , \ci_a[22] , 
        \ci_a[21] , \ci_a[20] , \ci_a[19] , \ci_a[18] , \ci_a[17] , \ci_a[16] , 
        \ci_a[15] , \ci_a[14] , \ci_a[13] , \ci_a[12] , \ci_a[11] , \ci_a[10] , 
        \ci_a[9] , \ci_a[8] , \ci_a[7] , \ci_a[6] , \ci_a[5] , \ci_a[4] , 
        \ci_a[3] , \ci_a[2] , \ci_a[1] , \ci_a[0] , \ci_wd[63] , \ci_wd[62] , 
        \ci_wd[61] , \ci_wd[60] , \ci_wd[59] , \ci_wd[58] , \ci_wd[57] , 
        \ci_wd[56] , \ci_wd[55] , \ci_wd[54] , \ci_wd[53] , \ci_wd[52] , 
        \ci_wd[51] , \ci_wd[50] , \ci_wd[49] , \ci_wd[48] , \ci_wd[47] , 
        \ci_wd[46] , \ci_wd[45] , \ci_wd[44] , \ci_wd[43] , \ci_wd[42] , 
        \ci_wd[41] , \ci_wd[40] , \ci_wd[39] , \ci_wd[38] , \ci_wd[37] , 
        \ci_wd[36] , \ci_wd[35] , \ci_wd[34] , \ci_wd[33] , \ci_wd[32] , 
        \ci_wd[31] , \ci_wd[30] , \ci_wd[29] , \ci_wd[28] , \ci_wd[27] , 
        \ci_wd[26] , \ci_wd[25] , \ci_wd[24] , \ci_wd[23] , \ci_wd[22] , 
        \ci_wd[21] , \ci_wd[20] , \ci_wd[19] , \ci_wd[18] , \ci_wd[17] , 
        \ci_wd[16] , \ci_wd[15] , \ci_wd[14] , \ci_wd[13] , \ci_wd[12] , 
        \ci_wd[11] , \ci_wd[10] , \ci_wd[9] , \ci_wd[8] , \ci_wd[7] , 
        \ci_wd[6] , \ci_wd[5] , \ci_wd[4] , \ci_wd[3] , \ci_wd[2] , \ci_wd[1] , 
        \ci_wd[0] , \ci_pred[1] , \ci_pred[0] , \ci_col[5] , \ci_col[4] , 
        \ci_col[3] , \ci_col[2] , \ci_col[1] , \ci_col[0] , ci_ack, 
        \ri_err[1] , \ri_err[0] , \ri_rnw[1] , \ri_rnw[0] , \ri_rd[63] , 
        \ri_rd[62] , \ri_rd[61] , \ri_rd[60] , \ri_rd[59] , \ri_rd[58] , 
        \ri_rd[57] , \ri_rd[56] , \ri_rd[55] , \ri_rd[54] , \ri_rd[53] , 
        \ri_rd[52] , \ri_rd[51] , \ri_rd[50] , \ri_rd[49] , \ri_rd[48] , 
        \ri_rd[47] , \ri_rd[46] , \ri_rd[45] , \ri_rd[44] , \ri_rd[43] , 
        \ri_rd[42] , \ri_rd[41] , \ri_rd[40] , \ri_rd[39] , \ri_rd[38] , 
        \ri_rd[37] , \ri_rd[36] , \ri_rd[35] , \ri_rd[34] , \ri_rd[33] , 
        \ri_rd[32] , \ri_rd[31] , \ri_rd[30] , \ri_rd[29] , \ri_rd[28] , 
        \ri_rd[27] , \ri_rd[26] , \ri_rd[25] , \ri_rd[24] , \ri_rd[23] , 
        \ri_rd[22] , \ri_rd[21] , \ri_rd[20] , \ri_rd[19] , \ri_rd[18] , 
        \ri_rd[17] , \ri_rd[16] , \ri_rd[15] , \ri_rd[14] , \ri_rd[13] , 
        \ri_rd[12] , \ri_rd[11] , \ri_rd[10] , \ri_rd[9] , \ri_rd[8] , 
        \ri_rd[7] , \ri_rd[6] , \ri_rd[5] , \ri_rd[4] , \ri_rd[3] , \ri_rd[2] , 
        \ri_rd[1] , \ri_rd[0] , ri_ack, reset, nroute_ack, routetx_req, 
        routetx_ack, \route[4] , \route[1] , \route[0] , \i_eh[2] , \i_eh[1] , 
        \i_eh[0] , \i_el[3] , \i_el[2] , \i_el[1] , \i_el[0] , \i_rh[3] , 
        \i_rh[2] , \i_rh[1] , \i_rl[3] , \i_rl[2] , \i_rl[1] , \i_rl[0] ;
    wire SYNOPSYS_UNCONNECTED_1 , SYNOPSYS_UNCONNECTED_2 , 
	SYNOPSYS_UNCONNECTED_3 , SYNOPSYS_UNCONNECTED_4 ;
    assign mr_rty = 1'b0;
    assign mr_acc = 1'b0;
    assign mr_ts[2] = 1'b0;
    assign mr_ts[1] = 1'b0;
    assign mr_ts[0] = 1'b0;
    assign mr_sel[3] = 1'b0;
    assign mr_sel[2] = 1'b0;
    assign mr_sel[1] = 1'b0;
    assign mr_sel[0] = 1'b0;
    inv_2 U1 ( .x(reset), .a(nReset) );
    m2cp_iport master2chainif ( .req_in(mc_req), .ts_o(mc_ts), .sel_o(mc_sel), 
        .mult_o(mc_mult), .we_o(mc_we), .prd_o(mc_prd), .seq_o(mc_seq), 
        .adr_o(mc_adr), .dat_o(mc_dat), .ain(mc_ack), .ic_seq({\ci_seq[1] , 
        \ci_seq[0] }), .ic_pred({\ci_pred[1] , \ci_pred[0] }), .ic_size({
        \ci_size[3] , \ci_size[2] , \ci_size[1] , \ci_size[0] }), .ic_itag({
        \ci_itag[9] , \ci_itag[8] , \ci_itag[7] , \ci_itag[6] , \ci_itag[5] , 
        \ci_itag[4] , \ci_itag[3] , \ci_itag[2] , \ci_itag[1] , \ci_itag[0] }), 
        .ic_wd({\ci_wd[63] , \ci_wd[62] , \ci_wd[61] , \ci_wd[60] , 
        \ci_wd[59] , \ci_wd[58] , \ci_wd[57] , \ci_wd[56] , \ci_wd[55] , 
        \ci_wd[54] , \ci_wd[53] , \ci_wd[52] , \ci_wd[51] , \ci_wd[50] , 
        \ci_wd[49] , \ci_wd[48] , \ci_wd[47] , \ci_wd[46] , \ci_wd[45] , 
        \ci_wd[44] , \ci_wd[43] , \ci_wd[42] , \ci_wd[41] , \ci_wd[40] , 
        \ci_wd[39] , \ci_wd[38] , \ci_wd[37] , \ci_wd[36] , \ci_wd[35] , 
        \ci_wd[34] , \ci_wd[33] , \ci_wd[32] , \ci_wd[31] , \ci_wd[30] , 
        \ci_wd[29] , \ci_wd[28] , \ci_wd[27] , \ci_wd[26] , \ci_wd[25] , 
        \ci_wd[24] , \ci_wd[23] , \ci_wd[22] , \ci_wd[21] , \ci_wd[20] , 
        \ci_wd[19] , \ci_wd[18] , \ci_wd[17] , \ci_wd[16] , \ci_wd[15] , 
        \ci_wd[14] , \ci_wd[13] , \ci_wd[12] , \ci_wd[11] , \ci_wd[10] , 
        \ci_wd[9] , \ci_wd[8] , \ci_wd[7] , \ci_wd[6] , \ci_wd[5] , \ci_wd[4] , 
        \ci_wd[3] , \ci_wd[2] , \ci_wd[1] , \ci_wd[0] }), .ic_lock({
        \ci_lock[1] , \ci_lock[0] }), .ic_a({\ci_a[63] , \ci_a[62] , 
        \ci_a[61] , \ci_a[60] , \ci_a[59] , \ci_a[58] , \ci_a[57] , \ci_a[56] , 
        \ci_a[55] , \ci_a[54] , \ci_a[53] , \ci_a[52] , \ci_a[51] , \ci_a[50] , 
        \ci_a[49] , \ci_a[48] , \ci_a[47] , \ci_a[46] , \ci_a[45] , \ci_a[44] , 
        \ci_a[43] , \ci_a[42] , \ci_a[41] , \ci_a[40] , \ci_a[39] , \ci_a[38] , 
        \ci_a[37] , \ci_a[36] , \ci_a[35] , \ci_a[34] , \ci_a[33] , \ci_a[32] , 
        \ci_a[31] , \ci_a[30] , \ci_a[29] , \ci_a[28] , \ci_a[27] , \ci_a[26] , 
        \ci_a[25] , \ci_a[24] , \ci_a[23] , \ci_a[22] , \ci_a[21] , \ci_a[20] , 
        \ci_a[19] , \ci_a[18] , \ci_a[17] , \ci_a[16] , \ci_a[15] , \ci_a[14] , 
        \ci_a[13] , \ci_a[12] , \ci_a[11] , \ci_a[10] , \ci_a[9] , \ci_a[8] , 
        \ci_a[7] , \ci_a[6] , \ci_a[5] , \ci_a[4] , \ci_a[3] , \ci_a[2] , 
        \ci_a[1] , \ci_a[0] }), .ic_rnw({\ci_rnw[1] , \ci_rnw[0] }), .ic_col({
        \ci_col[5] , \ci_col[4] , \ci_col[3] , \ci_col[2] , \ci_col[1] , 
        \ci_col[0] }), .ic_ack(ci_ack), .req_out(mr_req), .we_i(mr_we), 
        .err_i(mr_err), .dat_i(mr_dat), .aout(mr_ack), .ir_rd({\ri_rd[63] , 
        \ri_rd[62] , \ri_rd[61] , \ri_rd[60] , \ri_rd[59] , \ri_rd[58] , 
        \ri_rd[57] , \ri_rd[56] , \ri_rd[55] , \ri_rd[54] , \ri_rd[53] , 
        \ri_rd[52] , \ri_rd[51] , \ri_rd[50] , \ri_rd[49] , \ri_rd[48] , 
        \ri_rd[47] , \ri_rd[46] , \ri_rd[45] , \ri_rd[44] , \ri_rd[43] , 
        \ri_rd[42] , \ri_rd[41] , \ri_rd[40] , \ri_rd[39] , \ri_rd[38] , 
        \ri_rd[37] , \ri_rd[36] , \ri_rd[35] , \ri_rd[34] , \ri_rd[33] , 
        \ri_rd[32] , \ri_rd[31] , \ri_rd[30] , \ri_rd[29] , \ri_rd[28] , 
        \ri_rd[27] , \ri_rd[26] , \ri_rd[25] , \ri_rd[24] , \ri_rd[23] , 
        \ri_rd[22] , \ri_rd[21] , \ri_rd[20] , \ri_rd[19] , \ri_rd[18] , 
        \ri_rd[17] , \ri_rd[16] , \ri_rd[15] , \ri_rd[14] , \ri_rd[13] , 
        \ri_rd[12] , \ri_rd[11] , \ri_rd[10] , \ri_rd[9] , \ri_rd[8] , 
        \ri_rd[7] , \ri_rd[6] , \ri_rd[5] , \ri_rd[4] , \ri_rd[3] , \ri_rd[2] , 
        \ri_rd[1] , \ri_rd[0] }), .ir_err({\ri_err[1] , \ri_err[0] }), 
        .ir_rnw({\ri_rnw[1] , \ri_rnw[0] }), .ir_ack(ri_ack), .tag_id(tag_id), 
        .reset(reset) );
    i_adec_iport dec ( .e_h({SYNOPSYS_UNCONNECTED_1, \i_eh[2] , \i_eh[1] , 
        \i_eh[0] }), .e_l({\i_el[3] , \i_el[2] , \i_el[1] , \i_el[0] }), .r_h(
        {\i_rh[3] , \i_rh[2] , \i_rh[1] , SYNOPSYS_UNCONNECTED_2}), .r_l({
        \i_rl[3] , \i_rl[2] , \i_rl[1] , \i_rl[0] }), .ah({\ci_a[63] , 
        \ci_a[62] , \ci_a[61] , \ci_a[60] , \ci_a[59] , \ci_a[58] , \ci_a[57] , 
        \ci_a[56] , \ci_a[55] , \ci_a[54] , \ci_a[53] , \ci_a[52] , \ci_a[51] , 
        \ci_a[50] , \ci_a[49] , \ci_a[48] , \ci_a[47] , \ci_a[46] , \ci_a[45] , 
        \ci_a[44] , \ci_a[43] , \ci_a[42] , \ci_a[41] , \ci_a[40] , \ci_a[39] , 
        \ci_a[38] , \ci_a[37] , \ci_a[36] , \ci_a[35] , \ci_a[34] , \ci_a[33] , 
        \ci_a[32] }), .al({\ci_a[31] , \ci_a[30] , \ci_a[29] , \ci_a[28] , 
        \ci_a[27] , \ci_a[26] , \ci_a[25] , \ci_a[24] , \ci_a[23] , \ci_a[22] , 
        \ci_a[21] , \ci_a[20] , \ci_a[19] , \ci_a[18] , \ci_a[17] , \ci_a[16] , 
        \ci_a[15] , \ci_a[14] , \ci_a[13] , \ci_a[12] , \ci_a[11] , \ci_a[10] , 
        \ci_a[9] , \ci_a[8] , \ci_a[7] , \ci_a[6] , \ci_a[5] , \ci_a[4] , 
        \ci_a[3] , \ci_a[2] , \ci_a[1] , \ci_a[0] }), .e_bare(e_bare), .e_dm(
        e_dm), .e_im(e_im), .e_wish(e_wish), .r_bare(r_bare), .r_dm(r_dm), 
        .r_im(r_im), .r_wish(r_wish), .force_bare(force_bare) );
    route_tx_iport rt ( .o({\route[4] , SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, \route[1] , \route[0] }), .rtxack(routetx_ack), 
        .e_h({1'b0, \i_eh[2] , \i_eh[1] , \i_eh[0] }), .e_l({\i_el[3] , 
        \i_el[2] , \i_el[1] , \i_el[0] }), .noa(nroute_ack), .r_h({\i_rh[3] , 
        \i_rh[2] , \i_rh[1] , 1'b0}), .r_l({\i_rl[3] , \i_rl[2] , \i_rl[1] , 
        \i_rl[0] }), .rtxreq(routetx_req) );
    initiator_iport it ( .cack(ci_ack), .chaincommand(chaincommand), .err({
        \ri_err[1] , \ri_err[0] }), .nchainresponseack(nchainresponseack), 
        .nrouteack(nroute_ack), .rd({\ri_rd[63] , \ri_rd[62] , \ri_rd[61] , 
        \ri_rd[60] , \ri_rd[59] , \ri_rd[58] , \ri_rd[57] , \ri_rd[56] , 
        \ri_rd[55] , \ri_rd[54] , \ri_rd[53] , \ri_rd[52] , \ri_rd[51] , 
        \ri_rd[50] , \ri_rd[49] , \ri_rd[48] , \ri_rd[47] , \ri_rd[46] , 
        \ri_rd[45] , \ri_rd[44] , \ri_rd[43] , \ri_rd[42] , \ri_rd[41] , 
        \ri_rd[40] , \ri_rd[39] , \ri_rd[38] , \ri_rd[37] , \ri_rd[36] , 
        \ri_rd[35] , \ri_rd[34] , \ri_rd[33] , \ri_rd[32] , \ri_rd[31] , 
        \ri_rd[30] , \ri_rd[29] , \ri_rd[28] , \ri_rd[27] , \ri_rd[26] , 
        \ri_rd[25] , \ri_rd[24] , \ri_rd[23] , \ri_rd[22] , \ri_rd[21] , 
        \ri_rd[20] , \ri_rd[19] , \ri_rd[18] , \ri_rd[17] , \ri_rd[16] , 
        \ri_rd[15] , \ri_rd[14] , \ri_rd[13] , \ri_rd[12] , \ri_rd[11] , 
        \ri_rd[10] , \ri_rd[9] , \ri_rd[8] , \ri_rd[7] , \ri_rd[6] , 
        \ri_rd[5] , \ri_rd[4] , \ri_rd[3] , \ri_rd[2] , \ri_rd[1] , \ri_rd[0] 
        }), .routetxreq(routetx_req), .rrnw({\ri_rnw[1] , \ri_rnw[0] }), .a({
        \ci_a[63] , \ci_a[62] , \ci_a[61] , \ci_a[60] , \ci_a[59] , \ci_a[58] , 
        \ci_a[57] , \ci_a[56] , \ci_a[55] , \ci_a[54] , \ci_a[53] , \ci_a[52] , 
        \ci_a[51] , \ci_a[50] , \ci_a[49] , \ci_a[48] , \ci_a[47] , \ci_a[46] , 
        \ci_a[45] , \ci_a[44] , \ci_a[43] , \ci_a[42] , \ci_a[41] , \ci_a[40] , 
        \ci_a[39] , \ci_a[38] , \ci_a[37] , \ci_a[36] , \ci_a[35] , \ci_a[34] , 
        \ci_a[33] , \ci_a[32] , \ci_a[31] , \ci_a[30] , \ci_a[29] , \ci_a[28] , 
        \ci_a[27] , \ci_a[26] , \ci_a[25] , \ci_a[24] , \ci_a[23] , \ci_a[22] , 
        \ci_a[21] , \ci_a[20] , \ci_a[19] , \ci_a[18] , \ci_a[17] , \ci_a[16] , 
        \ci_a[15] , \ci_a[14] , \ci_a[13] , \ci_a[12] , \ci_a[11] , \ci_a[10] , 
        \ci_a[9] , \ci_a[8] , \ci_a[7] , \ci_a[6] , \ci_a[5] , \ci_a[4] , 
        \ci_a[3] , \ci_a[2] , \ci_a[1] , \ci_a[0] }), .chainresponse(
        chainresponse), .col({\ci_col[5] , \ci_col[4] , \ci_col[3] , 
        \ci_col[2] , \ci_col[1] , \ci_col[0] }), .crnw({\ci_rnw[1] , 
        \ci_rnw[0] }), .itag({\ci_itag[9] , \ci_itag[8] , \ci_itag[7] , 
        \ci_itag[6] , \ci_itag[5] , \ci_itag[4] , \ci_itag[3] , \ci_itag[2] , 
        \ci_itag[1] , \ci_itag[0] }), .lock({\ci_lock[1] , \ci_lock[0] }), 
        .nReset(nReset), .nchaincommandack(nchaincommandack), .pred({
        \ci_pred[1] , \ci_pred[0] }), .rack(ri_ack), .route({\route[4] , 1'b0, 
        1'b0, \route[1] , \route[0] }), .routetxack(routetx_ack), .seq({
        \ci_seq[1] , \ci_seq[0] }), .size({\ci_size[3] , \ci_size[2] , 
        \ci_size[1] , \ci_size[0] }), .wd({\ci_wd[63] , \ci_wd[62] , 
        \ci_wd[61] , \ci_wd[60] , \ci_wd[59] , \ci_wd[58] , \ci_wd[57] , 
        \ci_wd[56] , \ci_wd[55] , \ci_wd[54] , \ci_wd[53] , \ci_wd[52] , 
        \ci_wd[51] , \ci_wd[50] , \ci_wd[49] , \ci_wd[48] , \ci_wd[47] , 
        \ci_wd[46] , \ci_wd[45] , \ci_wd[44] , \ci_wd[43] , \ci_wd[42] , 
        \ci_wd[41] , \ci_wd[40] , \ci_wd[39] , \ci_wd[38] , \ci_wd[37] , 
        \ci_wd[36] , \ci_wd[35] , \ci_wd[34] , \ci_wd[33] , \ci_wd[32] , 
        \ci_wd[31] , \ci_wd[30] , \ci_wd[29] , \ci_wd[28] , \ci_wd[27] , 
        \ci_wd[26] , \ci_wd[25] , \ci_wd[24] , \ci_wd[23] , \ci_wd[22] , 
        \ci_wd[21] , \ci_wd[20] , \ci_wd[19] , \ci_wd[18] , \ci_wd[17] , 
        \ci_wd[16] , \ci_wd[15] , \ci_wd[14] , \ci_wd[13] , \ci_wd[12] , 
        \ci_wd[11] , \ci_wd[10] , \ci_wd[9] , \ci_wd[8] , \ci_wd[7] , 
        \ci_wd[6] , \ci_wd[5] , \ci_wd[4] , \ci_wd[3] , \ci_wd[2] , \ci_wd[1] , 
        \ci_wd[0] }) );
endmodule


module i_adec_dport ( e_h, e_l, r_h, r_l, ah, al, e_bare, e_dm, e_im, e_wish, 
    r_bare, r_dm, r_im, r_wish, force_bare );
output [3:0] e_h;
output [3:0] e_l;
output [3:0] r_h;
output [3:0] r_l;
input  [31:0] ah;
input  [31:0] al;
input  [3:0] e_bare;
input  [3:0] e_dm;
input  [3:0] e_im;
input  [3:0] e_wish;
input  [3:0] r_bare;
input  [3:0] r_dm;
input  [3:0] r_im;
input  [3:0] r_wish;
input  force_bare;
    wire \e_l[2] , \e_h[0] , n12, \r_l[3] , \r_l[2] , \r_l[0] , im_i, dm_i, 
        wish_i, bare_i, n1, n2, n3, n6, n7, \e_l[3] , \e_l[0] , \e_h[2] ;
    assign e_h[3] = 1'b0;
    assign e_h[2] = \e_h[2] ;
    assign e_h[0] = \e_h[0] ;
    assign e_l[3] = \e_l[3] ;
    assign e_l[2] = \e_l[2] ;
    assign e_l[0] = \e_l[0] ;
    assign r_h[3] = \e_l[2] ;
    assign r_h[2] = \e_h[0] ;
    assign r_h[0] = 1'b0;
    assign r_l[3] = \e_h[2] ;
    assign r_l[2] = \e_l[0] ;
    assign r_l[0] = \e_l[3] ;
    ao222_1 \U1632/U18/U1/U1  ( .x(wish_i), .a(n6), .b(al[30]), .c(n6), .d(
        wish_i), .e(al[30]), .f(wish_i) );
    ao222_1 \U1633/U18/U1/U1  ( .x(bare_i), .a(n6), .b(ah[30]), .c(n6), .d(
        bare_i), .e(ah[30]), .f(bare_i) );
    ao222_1 \U1634/U18/U1/U1  ( .x(im_i), .a(al[11]), .b(n7), .c(al[11]), .d(
        im_i), .e(n7), .f(im_i) );
    ao222_1 \U1635/U18/U1/U1  ( .x(dm_i), .a(ah[11]), .b(n7), .c(ah[11]), .d(
        dm_i), .e(n7), .f(dm_i) );
    or3_1 U1 ( .x(\r_l[2] ), .a(wish_i), .b(bare_i), .c(force_bare) );
    or2_1 U2 ( .x(r_l[1]), .a(\e_l[0] ), .b(im_i) );
    or2_1 U3 ( .x(\r_l[0] ), .a(dm_i), .b(r_l[1]) );
    nor2_0 U4 ( .x(n1), .a(bare_i), .b(force_bare) );
    aoi21_1 U6 ( .x(n2), .a(n3), .b(im_i), .c(r_h[1]) );
    inv_0 U8 ( .x(n3), .a(force_bare) );
    nor2i_0 U9 ( .x(\r_l[3] ), .a(wish_i), .b(force_bare) );
    nor2i_0 U10 ( .x(n12), .a(dm_i), .b(force_bare) );
    inv_0 U11 ( .x(e_h[1]), .a(n1) );
    buf_1 U15 ( .x(n6), .a(ah[31]) );
    buf_1 U16 ( .x(n7), .a(al[31]) );
    nand2_2 U17 ( .x(\e_l[2] ), .a(n2), .b(n1) );
    buf_1 U18 ( .x(r_h[1]), .a(n12) );
    inv_2 U19 ( .x(\e_h[0] ), .a(n2) );
    buf_3 U20 ( .x(\e_l[3] ), .a(\r_l[0] ) );
    buf_3 U21 ( .x(\e_l[0] ), .a(\r_l[2] ) );
    buf_3 U22 ( .x(\e_h[2] ), .a(\r_l[3] ) );
    nand2i_2 U23 ( .x(e_l[1]), .a(\e_h[2] ), .b(n2) );
endmodule


module chain_selement_ga_8 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_4 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[1] , \c[0] ;
    chain_selement_ga_8 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_9 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_5 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[1] , \c[0] ;
    chain_selement_ga_9 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_10 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_6 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[1] , \c[0] ;
    chain_selement_ga_10 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_11 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_7 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[1] , \c[0] ;
    chain_selement_ga_11 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_78 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_tx_dport ( o, rtxack, e_h, e_l, noa, r_h, r_l, rtxreq );
output [4:0] o;
input  [3:0] e_h;
input  [3:0] e_l;
input  [3:0] r_h;
input  [3:0] r_l;
input  noa, rtxreq;
output rtxack;
    wire \net52[0] , \net52[1] , \net55[0] , \net55[1] , \r3[2] , \r3[1] , 
        \r3[0] , \r0[2] , \r0[1] , \r0[0] , \r2[2] , \r2[1] , \r2[0] , 
        \last[0] , \last[1] , \last[2] , \last[3] , \last[4] , \r1[2] , 
        \r1[1] , \r1[0] , net6, eopsym, net9, net11, net16, net33, net60, 
        net40, net47, net50, \I8/nb , \I8/na , \I11/nc , \I11/nb , \I11/na , 
        \I7_0_/U25/U1/clr , \I7_0_/U25/U1/ob , \I7_1_/U25/U1/clr , 
        \I7_1_/U25/U1/ob ;
    assign o[3] = 1'b0;
    assign o[2] = 1'b0;
    route_symbol_4 I0 ( .o({\r3[2] , \r3[1] , \r3[0] }), .txack(net33), 
        .txack_last(\last[4] ), .e({e_h[3], e_l[3]}), .oa(net60), .r({r_h[3], 
        r_l[3]}), .txreq(rtxreq) );
    route_symbol_5 I1 ( .o({\r2[2] , \r2[1] , \r2[0] }), .txack(net40), 
        .txack_last(\last[3] ), .e({e_h[2], e_l[2]}), .oa(net60), .r({r_h[2], 
        r_l[2]}), .txreq(net33) );
    route_symbol_6 I2 ( .o({\r1[2] , \r1[1] , \r1[0] }), .txack(net47), 
        .txack_last(\last[2] ), .e({e_h[1], e_l[1]}), .oa(net60), .r({r_h[1], 
        r_l[1]}), .txreq(net40) );
    route_symbol_7 I3 ( .o({\r0[2] , \r0[1] , \r0[0] }), .txack(net50), 
        .txack_last(\last[1] ), .e({e_h[0], e_l[0]}), .oa(net60), .r({r_h[0], 
        r_l[0]}), .txreq(net47) );
    chain_selement_ga_78 I9 ( .Aa(\last[0] ), .Br(eopsym), .Ar(net50), .Ba(
        net60) );
    nor3_1 \I8/U27  ( .x(\I8/nb ), .a(o[4]), .b(o[3]), .c(o[2]) );
    nor2_1 \I8/U26  ( .x(\I8/na ), .a(o[1]), .b(o[0]) );
    nand2_2 \I8/U29  ( .x(net60), .a(\I8/nb ), .b(\I8/na ) );
    or2_1 \I13_0_/U12  ( .x(\net55[1] ), .a(\r1[0] ), .b(\r0[0] ) );
    or2_1 \I13_1_/U12  ( .x(\net55[0] ), .a(\r1[1] ), .b(\r0[1] ) );
    or2_1 \I14_0_/U12  ( .x(\net52[1] ), .a(\r3[0] ), .b(\r2[0] ) );
    or2_1 \I14_1_/U12  ( .x(\net52[0] ), .a(\r3[1] ), .b(\r2[1] ) );
    nand3_1 \I11/U31  ( .x(rtxack), .a(\I11/nc ), .b(\I11/nb ), .c(\I11/na )
         );
    inv_1 \I11/U33  ( .x(\I11/nc ), .a(\last[0] ) );
    nor2_1 \I11/U26  ( .x(\I11/na ), .a(\last[3] ), .b(\last[4] ) );
    nor2_1 \I11/U32  ( .x(\I11/nb ), .a(\last[1] ), .b(\last[2] ) );
    nor2_1 \I16/U5  ( .x(net16), .a(\r1[2] ), .b(\r0[2] ) );
    nor2_1 \I5/U5  ( .x(net11), .a(\r3[2] ), .b(\r2[2] ) );
    nand3_1 \I17/U9  ( .x(net9), .a(net6), .b(net11), .c(net16) );
    inv_1 \I18/U3  ( .x(net6), .a(eopsym) );
    oa31_1 \I7_0_/U25/U1/Uclr  ( .x(\I7_0_/U25/U1/clr ), .a(noa), .b(
        \net55[1] ), .c(\net52[1] ), .d(o[0]) );
    oaoi211_1 \I7_0_/U25/U1/Uaoi  ( .x(\I7_0_/U25/U1/ob ), .a(\net55[1] ), .b(
        \net52[1] ), .c(noa), .d(\I7_0_/U25/U1/clr ) );
    inv_2 \I7_0_/U25/U1/Ui  ( .x(o[0]), .a(\I7_0_/U25/U1/ob ) );
    oa31_1 \I7_1_/U25/U1/Uclr  ( .x(\I7_1_/U25/U1/clr ), .a(noa), .b(
        \net55[0] ), .c(\net52[0] ), .d(o[1]) );
    oaoi211_1 \I7_1_/U25/U1/Uaoi  ( .x(\I7_1_/U25/U1/ob ), .a(\net55[0] ), .b(
        \net52[0] ), .c(noa), .d(\I7_1_/U25/U1/clr ) );
    inv_2 \I7_1_/U25/U1/Ui  ( .x(o[1]), .a(\I7_1_/U25/U1/ob ) );
    ao222_1 \I15/U18/U1/U1  ( .x(o[4]), .a(noa), .b(net9), .c(noa), .d(o[4]), 
        .e(net9), .f(o[4]) );
endmodule


module chain_dr8bit_completion_24 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_25 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_26 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_27 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr32bit_completion_4 ( o, i );
input  [63:0] i;
output o;
    wire nx, \cd[3] , \cd[2] , ny, \cd[0] , \cd[1] , \U16/Z , \U6/Z , \U15/Z ;
    chain_dr8bit_completion_24 U11 ( .o(\cd[3] ), .i({i[63], i[62], i[61], 
        i[60], i[59], i[58], i[57], i[56], i[31], i[30], i[29], i[28], i[27], 
        i[26], i[25], i[24]}) );
    chain_dr8bit_completion_27 U14 ( .o(\cd[2] ), .i({i[55], i[54], i[53], 
        i[52], i[51], i[50], i[49], i[48], i[23], i[22], i[21], i[20], i[19], 
        i[18], i[17], i[16]}) );
    chain_dr8bit_completion_26 U13 ( .o(\cd[1] ), .i({i[47], i[46], i[45], 
        i[44], i[43], i[42], i[41], i[40], i[15], i[14], i[13], i[12], i[11], 
        i[10], i[9], i[8]}) );
    chain_dr8bit_completion_25 U12 ( .o(\cd[0] ), .i({i[39], i[38], i[37], 
        i[36], i[35], i[34], i[33], i[32], i[7], i[6], i[5], i[4], i[3], i[2], 
        i[1], i[0]}) );
    aoi222_1 \U16/U30/U1  ( .x(ny), .a(\cd[0] ), .b(\cd[1] ), .c(\cd[0] ), .d(
        \U16/Z ), .e(\cd[1] ), .f(\U16/Z ) );
    inv_1 \U16/U30/Uinv  ( .x(\U16/Z ), .a(ny) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(ny), .b(nx), .c(ny), .d(\U6/Z ), .e(nx), 
        .f(\U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U15/U30/U1  ( .x(nx), .a(\cd[3] ), .b(\cd[2] ), .c(\cd[3] ), .d(
        \U15/Z ), .e(\cd[2] ), .f(\U15/Z ) );
    inv_1 \U15/U30/Uinv  ( .x(\U15/Z ), .a(nx) );
endmodule


module chain_dr8bit_completion_28 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_29 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_30 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_31 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr32bit_completion_5 ( o, i );
input  [63:0] i;
output o;
    wire nx, \cd[3] , \cd[2] , ny, \cd[0] , \cd[1] , \U16/Z , \U6/Z , \U15/Z ;
    chain_dr8bit_completion_28 U11 ( .o(\cd[3] ), .i({i[63], i[62], i[61], 
        i[60], i[59], i[58], i[57], i[56], i[31], i[30], i[29], i[28], i[27], 
        i[26], i[25], i[24]}) );
    chain_dr8bit_completion_31 U14 ( .o(\cd[2] ), .i({i[55], i[54], i[53], 
        i[52], i[51], i[50], i[49], i[48], i[23], i[22], i[21], i[20], i[19], 
        i[18], i[17], i[16]}) );
    chain_dr8bit_completion_30 U13 ( .o(\cd[1] ), .i({i[47], i[46], i[45], 
        i[44], i[43], i[42], i[41], i[40], i[15], i[14], i[13], i[12], i[11], 
        i[10], i[9], i[8]}) );
    chain_dr8bit_completion_29 U12 ( .o(\cd[0] ), .i({i[39], i[38], i[37], 
        i[36], i[35], i[34], i[33], i[32], i[7], i[6], i[5], i[4], i[3], i[2], 
        i[1], i[0]}) );
    aoi222_1 \U16/U30/U1  ( .x(ny), .a(\cd[0] ), .b(\cd[1] ), .c(\cd[0] ), .d(
        \U16/Z ), .e(\cd[1] ), .f(\U16/Z ) );
    inv_1 \U16/U30/Uinv  ( .x(\U16/Z ), .a(ny) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(ny), .b(nx), .c(ny), .d(\U6/Z ), .e(nx), 
        .f(\U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U15/U30/U1  ( .x(nx), .a(\cd[3] ), .b(\cd[2] ), .c(\cd[3] ), .d(
        \U15/Z ), .e(\cd[2] ), .f(\U15/Z ) );
    inv_1 \U15/U30/Uinv  ( .x(\U15/Z ), .a(nx) );
endmodule


module chain_dr8bit_completion_52 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_53 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_selement_ga_42 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_43 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_44 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_45 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_46 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_47 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_48 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_49 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_50 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_51 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_icmux_1 ( ack, chainh, chainl, sendack, addr, col, itag, lock, 
    nReset, nia, pred, rnw, sendreq, seq, size, wd );
output [7:0] chainh;
output [7:0] chainl;
input  [63:0] addr;
input  [5:0] col;
input  [9:0] itag;
input  [1:0] lock;
input  [1:0] pred;
input  [1:0] rnw;
input  [1:0] seq;
input  [3:0] size;
input  [63:0] wd;
input  nReset, nia, sendreq;
output ack, sendack;
    wire \net207[0] , \net207[1] , \net207[2] , \net207[3] , \net207[4] , 
        \net207[5] , \net207[6] , \net207[7] , \net207[8] , \net207[9] , 
        \net207[10] , \net207[11] , \net207[12] , \net207[13] , \net207[14] , 
        \net207[15] , \bs[0] , \bs[1] , \bs[2] , \bs[3] , \bs[4] , \bs[5] , 
        \bs[6] , \bs[7] , \bs[8] , \net231[0] , \net231[1] , \net231[2] , 
        \net231[3] , \net231[4] , \net231[5] , \net231[6] , \net231[7] , 
        \net231[8] , \net231[9] , \net231[10] , \net231[11] , \net231[12] , 
        \net231[13] , \net231[14] , \net231[15] , \hdr[4] , \net234[0] , 
        \net234[1] , \net234[2] , \net234[3] , \net234[4] , \net234[5] , 
        \net234[6] , \net234[7] , \net234[8] , \net234[9] , \net234[10] , 
        \net234[11] , \net234[12] , \net234[13] , \net234[14] , \net234[15] , 
        \net217[0] , \net217[1] , \net217[2] , \net217[3] , \net217[4] , 
        \net217[5] , \net217[6] , \net217[7] , \net217[8] , \net217[9] , 
        \net217[10] , \net217[11] , \net217[12] , \net217[13] , \net217[14] , 
        \net217[15] , \net246[0] , \net246[1] , \net246[2] , \net246[3] , 
        \net246[4] , \net246[5] , \net246[6] , \net246[7] , \net246[8] , 
        \net246[9] , \net246[10] , \net246[11] , \net246[12] , \net246[13] , 
        \net246[14] , \net246[15] , \net243[0] , \net243[1] , \net243[2] , 
        \net243[3] , \net243[4] , \net243[5] , \net243[6] , \net243[7] , 
        \net243[8] , \net243[9] , \net243[10] , \net243[11] , \net243[12] , 
        \net243[13] , \net243[14] , \net243[15] , \net240[0] , \net240[1] , 
        \net240[2] , \net240[3] , \net240[4] , \net240[5] , \net240[6] , 
        \net240[7] , \net240[8] , \net240[9] , \net240[10] , \net240[11] , 
        \net240[12] , \net240[13] , \net240[14] , \net240[15] , \net219[0] , 
        \net219[1] , \net219[2] , \net219[3] , \net219[4] , \net219[5] , 
        \net219[6] , \net219[7] , \net219[8] , \net219[9] , \net219[10] , 
        \net219[11] , \net219[12] , \net219[13] , \net219[14] , \net219[15] , 
        \net237[0] , \net237[1] , \net237[2] , \net237[5] , \net237[6] , 
        \net237[7] , \net237[8] , \net237[9] , \net237[10] , \net237[11] , 
        \net237[12] , \net237[13] , \net237[14] , \net237[15] , \net222[0] , 
        \net222[1] , \net222[2] , \net222[3] , \net222[4] , \net222[5] , 
        \net222[6] , \net222[7] , \net222[8] , \net222[9] , \net222[10] , 
        \net222[11] , \net222[12] , \net222[13] , \net222[14] , \net222[15] , 
        \net225[0] , \net225[1] , \net225[2] , \net225[3] , \net225[4] , 
        \net225[5] , \net225[6] , \net225[7] , \net225[8] , \net225[9] , 
        \net225[10] , \net225[11] , \net225[12] , \net225[13] , \net225[14] , 
        \net225[15] , \net228[0] , \net228[1] , \net228[2] , \net228[3] , 
        \net228[4] , \net228[5] , \net228[6] , \net228[7] , \net228[8] , 
        \net228[9] , \net228[10] , \net228[11] , \net228[12] , \net228[13] , 
        \net228[14] , \net228[15] , \net212[0] , \net212[1] , \net212[2] , 
        \net212[3] , \net212[4] , \net212[5] , \net212[6] , \net212[7] , 
        \net212[8] , \net212[9] , \net212[10] , \net212[11] , \net212[12] , 
        \net212[13] , \net212[14] , \net212[15] , net138, net198, net176, 
        net132, net131, net136, net185, net187, net191, net293, net152, net146, 
        net148, net156, net160, net168, net172, net164, net289, net180, net189, 
        net249, net261, net251, net255, net253, net259, net269, net267, net263, 
        net265, \U40_0_/n5 , \U40_0_/n3 , \U40_0_/n4 , \U40_1_/n5 , 
        \U40_1_/n3 , \U40_1_/n4 , \U40_2_/n5 , \U40_2_/n3 , \U40_2_/n4 , 
        \U40_3_/n5 , \U40_3_/n3 , \U40_3_/n4 , \U40_4_/n5 , \U40_4_/n3 , 
        \U40_4_/n4 , \U40_5_/n5 , \U40_5_/n3 , \U40_5_/n4 , \U40_6_/n5 , 
        \U40_6_/n3 , \U40_6_/n4 , \U40_7_/n5 , \U40_7_/n3 , \U40_7_/n4 , 
        \U40_8_/n5 , \U40_8_/n3 , \U40_8_/n4 , \U40_9_/n5 , \U40_9_/n3 , 
        \U40_9_/n4 , \U40_10_/n5 , \U40_10_/n3 , \U40_10_/n4 , \U40_11_/n5 , 
        \U40_11_/n3 , \U40_11_/n4 , \U40_12_/n5 , \U40_12_/n3 , \U40_12_/n4 , 
        \U40_13_/n5 , \U40_13_/n3 , \U40_13_/n4 , \U40_14_/n5 , \U40_14_/n3 , 
        \U40_14_/n4 , \U40_15_/n5 , \U40_15_/n3 , \U40_15_/n4 , \U14_0_/n5 , 
        \U14_0_/n1 , \U14_0_/n2 , \U14_0_/n3 , \U14_0_/n4 , \U14_1_/n5 , 
        \U14_1_/n1 , \U14_1_/n2 , \U14_1_/n3 , \U14_1_/n4 , \U14_2_/n5 , 
        \U14_2_/n1 , \U14_2_/n2 , \U14_2_/n3 , \U14_2_/n4 , \U14_3_/n5 , 
        \U14_3_/n1 , \U14_3_/n2 , \U14_3_/n3 , \U14_3_/n4 , \U14_4_/n5 , 
        \U14_4_/n1 , \U14_4_/n2 , \U14_4_/n3 , \U14_4_/n4 , \U14_5_/n5 , 
        \U14_5_/n1 , \U14_5_/n2 , \U14_5_/n3 , \U14_5_/n4 , \U14_6_/n5 , 
        \U14_6_/n1 , \U14_6_/n2 , \U14_6_/n3 , \U14_6_/n4 , \U14_7_/n5 , 
        \U14_7_/n1 , \U14_7_/n2 , \U14_7_/n3 , \U14_7_/n4 , \U14_8_/n5 , 
        \U14_8_/n1 , \U14_8_/n2 , \U14_8_/n3 , \U14_8_/n4 , \U14_9_/n5 , 
        \U14_9_/n1 , \U14_9_/n2 , \U14_9_/n3 , \U14_9_/n4 , \U14_10_/n5 , 
        \U14_10_/n1 , \U14_10_/n2 , \U14_10_/n3 , \U14_10_/n4 , \U14_11_/n5 , 
        \U14_11_/n1 , \U14_11_/n2 , \U14_11_/n4 , \U14_12_/n5 , \U14_12_/n1 , 
        \U14_12_/n2 , \U14_12_/n4 , \U14_13_/n5 , \U14_13_/n1 , \U14_13_/n2 , 
        \U14_13_/n3 , \U14_13_/n4 , \U14_14_/n5 , \U14_14_/n1 , \U14_14_/n2 , 
        \U14_14_/n3 , \U14_14_/n4 , \U14_15_/n5 , \U14_15_/n1 , \U14_15_/n2 , 
        \U14_15_/n3 , \U14_15_/n4 , \U91_0_/n5 , \U91_0_/n1 , \U91_0_/n2 , 
        \U91_0_/n3 , \U91_0_/n4 , \U91_1_/n5 , \U91_1_/n1 , \U91_1_/n2 , 
        \U91_1_/n3 , \U91_1_/n4 , \U91_2_/n5 , \U91_2_/n1 , \U91_2_/n2 , 
        \U91_2_/n3 , \U91_2_/n4 , \U91_3_/n5 , \U91_3_/n1 , \U91_3_/n2 , 
        \U91_3_/n3 , \U91_3_/n4 , \U91_4_/n5 , \U91_4_/n1 , \U91_4_/n2 , 
        \U91_4_/n3 , \U91_4_/n4 , \U91_5_/n5 , \U91_5_/n1 , \U91_5_/n2 , 
        \U91_5_/n3 , \U91_5_/n4 , \U91_6_/n5 , \U91_6_/n1 , \U91_6_/n2 , 
        \U91_6_/n3 , \U91_6_/n4 , \U91_7_/n5 , \U91_7_/n1 , \U91_7_/n2 , 
        \U91_7_/n3 , \U91_7_/n4 , \U91_8_/n5 , \U91_8_/n1 , \U91_8_/n2 , 
        \U91_8_/n3 , \U91_8_/n4 , \U91_9_/n5 , \U91_9_/n1 , \U91_9_/n2 , 
        \U91_9_/n3 , \U91_9_/n4 , \U91_10_/n5 , \U91_10_/n1 , \U91_10_/n2 , 
        \U91_10_/n3 , \U91_10_/n4 , \U91_11_/n5 , \U91_11_/n1 , \U91_11_/n2 , 
        \U91_11_/n3 , \U91_11_/n4 , \U91_12_/n5 , \U91_12_/n1 , \U91_12_/n2 , 
        \U91_12_/n3 , \U91_12_/n4 , \U91_13_/n5 , \U91_13_/n1 , \U91_13_/n2 , 
        \U91_13_/n3 , \U91_13_/n4 , \U91_14_/n5 , \U91_14_/n1 , \U91_14_/n2 , 
        \U91_14_/n3 , \U91_14_/n4 , \U91_15_/n5 , \U91_15_/n1 , \U91_15_/n2 , 
        \U91_15_/n3 , \U91_15_/n4 , \U148/U21/nr , \U148/U21/nd , 
        \U148/U21/n2 , \U151/Z , n1;
    chain_selement_ga_43 U163 ( .Aa(net152), .Br(net146), .Ar(net148), .Ba(n1)
         );
    chain_selement_ga_44 U164 ( .Aa(net156), .Br(\bs[1] ), .Ar(net152), .Ba(
        net138) );
    chain_selement_ga_45 U165 ( .Aa(net160), .Br(\bs[2] ), .Ar(net156), .Ba(n1
        ) );
    chain_selement_ga_46 U166 ( .Aa(net168), .Br(\bs[3] ), .Ar(net160), .Ba(
        net138) );
    chain_selement_ga_50 U170 ( .Aa(net172), .Br(\bs[7] ), .Ar(net164), .Ba(
        net138) );
    chain_selement_ga_47 U167 ( .Aa(net132), .Br(\bs[4] ), .Ar(net168), .Ba(
        net138) );
    chain_selement_ga_51 U171 ( .Aa(net289), .Br(\bs[8] ), .Ar(net172), .Ba(
        net138) );
    chain_selement_ga_48 U168 ( .Aa(net180), .Br(\bs[5] ), .Ar(net176), .Ba(
        net138) );
    chain_selement_ga_49 U169 ( .Aa(net164), .Br(\bs[6] ), .Ar(net180), .Ba(n1
        ) );
    chain_selement_ga_42 U161 ( .Aa(net148), .Br(\bs[0] ), .Ar(\hdr[4] ), .Ba(
        n1) );
    chain_dr8bit_completion_52 U119 ( .o(net185), .i({col[5], col[4], col[3], 
        itag[9], itag[8], itag[7], itag[6], itag[5], col[2], col[1], col[0], 
        itag[4], itag[3], itag[2], itag[1], itag[0]}) );
    chain_dr8bit_completion_53 U147 ( .o(net187), .i({size[3], size[2], rnw[1], 
        1'b0, 1'b0, lock[1], pred[1], seq[1], size[1], size[0], rnw[0], 
        \hdr[4] , \hdr[4] , lock[0], pred[0], seq[0]}) );
    chain_dr32bit_completion_4 U117 ( .o(net189), .i(wd) );
    chain_dr32bit_completion_5 U118 ( .o(net191), .i(addr) );
    or2_4 \U122/U12  ( .x(net293), .a(net189), .b(net131) );
    or2_4 \U53/U12  ( .x(sendack), .a(net131), .b(net289) );
    and2_1 \U32_0_/U8  ( .x(\net246[15] ), .a(itag[0]), .b(net265) );
    and2_1 \U32_1_/U8  ( .x(\net246[14] ), .a(itag[1]), .b(net265) );
    and2_1 \U32_2_/U8  ( .x(\net246[13] ), .a(itag[2]), .b(net265) );
    and2_1 \U32_3_/U8  ( .x(\net246[12] ), .a(itag[3]), .b(net265) );
    and2_1 \U32_4_/U8  ( .x(\net246[11] ), .a(itag[4]), .b(net265) );
    and2_1 \U32_5_/U8  ( .x(\net246[10] ), .a(col[0]), .b(net265) );
    and2_1 \U32_6_/U8  ( .x(\net246[9] ), .a(col[1]), .b(net265) );
    and2_1 \U32_7_/U8  ( .x(\net246[8] ), .a(col[2]), .b(net265) );
    and2_1 \U32_8_/U8  ( .x(\net246[7] ), .a(itag[5]), .b(net265) );
    and2_1 \U32_9_/U8  ( .x(\net246[6] ), .a(itag[6]), .b(net265) );
    and2_1 \U32_10_/U8  ( .x(\net246[5] ), .a(itag[7]), .b(net265) );
    and2_1 \U32_11_/U8  ( .x(\net246[4] ), .a(itag[8]), .b(net265) );
    and2_1 \U32_12_/U8  ( .x(\net246[3] ), .a(itag[9]), .b(net265) );
    and2_1 \U32_13_/U8  ( .x(\net246[2] ), .a(col[3]), .b(net265) );
    and2_1 \U32_14_/U8  ( .x(\net246[1] ), .a(col[4]), .b(net265) );
    and2_1 \U32_15_/U8  ( .x(\net246[0] ), .a(col[5]), .b(net265) );
    and2_1 \U76_0_/U8  ( .x(\net243[15] ), .a(wd[8]), .b(net263) );
    and2_1 \U76_1_/U8  ( .x(\net243[14] ), .a(wd[9]), .b(net263) );
    and2_1 \U76_2_/U8  ( .x(\net243[13] ), .a(wd[10]), .b(net263) );
    and2_1 \U76_3_/U8  ( .x(\net243[12] ), .a(wd[11]), .b(net263) );
    and2_1 \U76_4_/U8  ( .x(\net243[11] ), .a(wd[12]), .b(net263) );
    and2_1 \U76_5_/U8  ( .x(\net243[10] ), .a(wd[13]), .b(net263) );
    and2_1 \U76_6_/U8  ( .x(\net243[9] ), .a(wd[14]), .b(net263) );
    and2_1 \U76_7_/U8  ( .x(\net243[8] ), .a(wd[15]), .b(net263) );
    and2_1 \U76_8_/U8  ( .x(\net243[7] ), .a(wd[40]), .b(net263) );
    and2_1 \U76_9_/U8  ( .x(\net243[6] ), .a(wd[41]), .b(net263) );
    and2_1 \U76_10_/U8  ( .x(\net243[5] ), .a(wd[42]), .b(net263) );
    and2_1 \U76_11_/U8  ( .x(\net243[4] ), .a(wd[43]), .b(net263) );
    and2_1 \U76_12_/U8  ( .x(\net243[3] ), .a(wd[44]), .b(net263) );
    and2_1 \U76_13_/U8  ( .x(\net243[2] ), .a(wd[45]), .b(net263) );
    and2_1 \U76_14_/U8  ( .x(\net243[1] ), .a(wd[46]), .b(net263) );
    and2_1 \U76_15_/U8  ( .x(\net243[0] ), .a(wd[47]), .b(net263) );
    and2_1 \U80_0_/U8  ( .x(\net240[15] ), .a(wd[16]), .b(net267) );
    and2_1 \U80_1_/U8  ( .x(\net240[14] ), .a(wd[17]), .b(net267) );
    and2_1 \U80_2_/U8  ( .x(\net240[13] ), .a(wd[18]), .b(net267) );
    and2_1 \U80_3_/U8  ( .x(\net240[12] ), .a(wd[19]), .b(net267) );
    and2_1 \U80_4_/U8  ( .x(\net240[11] ), .a(wd[20]), .b(net267) );
    and2_1 \U80_5_/U8  ( .x(\net240[10] ), .a(wd[21]), .b(net267) );
    and2_1 \U80_6_/U8  ( .x(\net240[9] ), .a(wd[22]), .b(net267) );
    and2_1 \U80_7_/U8  ( .x(\net240[8] ), .a(wd[23]), .b(net267) );
    and2_1 \U80_8_/U8  ( .x(\net240[7] ), .a(wd[48]), .b(net267) );
    and2_1 \U80_9_/U8  ( .x(\net240[6] ), .a(wd[49]), .b(net267) );
    and2_1 \U80_10_/U8  ( .x(\net240[5] ), .a(wd[50]), .b(net267) );
    and2_1 \U80_11_/U8  ( .x(\net240[4] ), .a(wd[51]), .b(net267) );
    and2_1 \U80_12_/U8  ( .x(\net240[3] ), .a(wd[52]), .b(net267) );
    and2_1 \U80_13_/U8  ( .x(\net240[2] ), .a(wd[53]), .b(net267) );
    and2_1 \U80_14_/U8  ( .x(\net240[1] ), .a(wd[54]), .b(net267) );
    and2_1 \U80_15_/U8  ( .x(\net240[0] ), .a(wd[55]), .b(net267) );
    and2_1 \U128_0_/U8  ( .x(\net237[15] ), .a(seq[0]), .b(net269) );
    and2_1 \U128_1_/U8  ( .x(\net237[14] ), .a(pred[0]), .b(net269) );
    and2_1 \U128_2_/U8  ( .x(\net237[13] ), .a(lock[0]), .b(net269) );
    and2_1 \U128_3_/U8  ( .x(\net237[12] ), .a(\hdr[4] ), .b(net269) );
    and2_1 \U128_4_/U8  ( .x(\net237[11] ), .a(\hdr[4] ), .b(net269) );
    and2_1 \U128_5_/U8  ( .x(\net237[10] ), .a(rnw[0]), .b(net269) );
    and2_1 \U128_6_/U8  ( .x(\net237[9] ), .a(size[0]), .b(net269) );
    and2_1 \U128_7_/U8  ( .x(\net237[8] ), .a(size[1]), .b(net269) );
    and2_1 \U128_8_/U8  ( .x(\net237[7] ), .a(seq[1]), .b(net269) );
    and2_1 \U128_9_/U8  ( .x(\net237[6] ), .a(pred[1]), .b(net269) );
    and2_1 \U128_10_/U8  ( .x(\net237[5] ), .a(lock[1]), .b(net269) );
    and2_1 \U128_13_/U8  ( .x(\net237[2] ), .a(rnw[1]), .b(net269) );
    and2_1 \U128_14_/U8  ( .x(\net237[1] ), .a(size[2]), .b(net269) );
    and2_1 \U128_15_/U8  ( .x(\net237[0] ), .a(size[3]), .b(net269) );
    and2_1 \U37_0_/U8  ( .x(\net234[15] ), .a(addr[8]), .b(net259) );
    and2_1 \U37_1_/U8  ( .x(\net234[14] ), .a(addr[9]), .b(net259) );
    and2_1 \U37_2_/U8  ( .x(\net234[13] ), .a(addr[10]), .b(net259) );
    and2_1 \U37_3_/U8  ( .x(\net234[12] ), .a(addr[11]), .b(net259) );
    and2_1 \U37_4_/U8  ( .x(\net234[11] ), .a(addr[12]), .b(net259) );
    and2_1 \U37_5_/U8  ( .x(\net234[10] ), .a(addr[13]), .b(net259) );
    and2_1 \U37_6_/U8  ( .x(\net234[9] ), .a(addr[14]), .b(net259) );
    and2_1 \U37_7_/U8  ( .x(\net234[8] ), .a(addr[15]), .b(net259) );
    and2_1 \U37_8_/U8  ( .x(\net234[7] ), .a(addr[40]), .b(net259) );
    and2_1 \U37_9_/U8  ( .x(\net234[6] ), .a(addr[41]), .b(net259) );
    and2_1 \U37_10_/U8  ( .x(\net234[5] ), .a(addr[42]), .b(net259) );
    and2_1 \U37_11_/U8  ( .x(\net234[4] ), .a(addr[43]), .b(net259) );
    and2_1 \U37_12_/U8  ( .x(\net234[3] ), .a(addr[44]), .b(net259) );
    and2_1 \U37_13_/U8  ( .x(\net234[2] ), .a(addr[45]), .b(net259) );
    and2_1 \U37_14_/U8  ( .x(\net234[1] ), .a(addr[46]), .b(net259) );
    and2_1 \U37_15_/U8  ( .x(\net234[0] ), .a(addr[47]), .b(net259) );
    and2_1 \U33_0_/U8  ( .x(\net231[15] ), .a(addr[16]), .b(net253) );
    and2_1 \U33_1_/U8  ( .x(\net231[14] ), .a(addr[17]), .b(net253) );
    and2_1 \U33_2_/U8  ( .x(\net231[13] ), .a(addr[18]), .b(net253) );
    and2_1 \U33_3_/U8  ( .x(\net231[12] ), .a(addr[19]), .b(net253) );
    and2_1 \U33_4_/U8  ( .x(\net231[11] ), .a(addr[20]), .b(net253) );
    and2_1 \U33_5_/U8  ( .x(\net231[10] ), .a(addr[21]), .b(net253) );
    and2_1 \U33_6_/U8  ( .x(\net231[9] ), .a(addr[22]), .b(net253) );
    and2_1 \U33_7_/U8  ( .x(\net231[8] ), .a(addr[23]), .b(net253) );
    and2_1 \U33_8_/U8  ( .x(\net231[7] ), .a(addr[48]), .b(net253) );
    and2_1 \U33_9_/U8  ( .x(\net231[6] ), .a(addr[49]), .b(net253) );
    and2_1 \U33_10_/U8  ( .x(\net231[5] ), .a(addr[50]), .b(net253) );
    and2_1 \U33_11_/U8  ( .x(\net231[4] ), .a(addr[51]), .b(net253) );
    and2_1 \U33_12_/U8  ( .x(\net231[3] ), .a(addr[52]), .b(net253) );
    and2_1 \U33_13_/U8  ( .x(\net231[2] ), .a(addr[53]), .b(net253) );
    and2_1 \U33_14_/U8  ( .x(\net231[1] ), .a(addr[54]), .b(net253) );
    and2_1 \U33_15_/U8  ( .x(\net231[0] ), .a(addr[55]), .b(net253) );
    and2_1 \U81_0_/U8  ( .x(\net228[15] ), .a(wd[24]), .b(net255) );
    and2_1 \U81_1_/U8  ( .x(\net228[14] ), .a(wd[25]), .b(net255) );
    and2_1 \U81_2_/U8  ( .x(\net228[13] ), .a(wd[26]), .b(net255) );
    and2_1 \U81_3_/U8  ( .x(\net228[12] ), .a(wd[27]), .b(net255) );
    and2_1 \U81_4_/U8  ( .x(\net228[11] ), .a(wd[28]), .b(net255) );
    and2_1 \U81_5_/U8  ( .x(\net228[10] ), .a(wd[29]), .b(net255) );
    and2_1 \U81_6_/U8  ( .x(\net228[9] ), .a(wd[30]), .b(net255) );
    and2_1 \U81_7_/U8  ( .x(\net228[8] ), .a(wd[31]), .b(net255) );
    and2_1 \U81_8_/U8  ( .x(\net228[7] ), .a(wd[56]), .b(net255) );
    and2_1 \U81_9_/U8  ( .x(\net228[6] ), .a(wd[57]), .b(net255) );
    and2_1 \U81_10_/U8  ( .x(\net228[5] ), .a(wd[58]), .b(net255) );
    and2_1 \U81_11_/U8  ( .x(\net228[4] ), .a(wd[59]), .b(net255) );
    and2_1 \U81_12_/U8  ( .x(\net228[3] ), .a(wd[60]), .b(net255) );
    and2_1 \U81_13_/U8  ( .x(\net228[2] ), .a(wd[61]), .b(net255) );
    and2_1 \U81_14_/U8  ( .x(\net228[1] ), .a(wd[62]), .b(net255) );
    and2_1 \U81_15_/U8  ( .x(\net228[0] ), .a(wd[63]), .b(net255) );
    and2_1 \U34_0_/U8  ( .x(\net225[15] ), .a(addr[0]), .b(net251) );
    and2_1 \U34_1_/U8  ( .x(\net225[14] ), .a(addr[1]), .b(net251) );
    and2_1 \U34_2_/U8  ( .x(\net225[13] ), .a(addr[2]), .b(net251) );
    and2_1 \U34_3_/U8  ( .x(\net225[12] ), .a(addr[3]), .b(net251) );
    and2_1 \U34_4_/U8  ( .x(\net225[11] ), .a(addr[4]), .b(net251) );
    and2_1 \U34_5_/U8  ( .x(\net225[10] ), .a(addr[5]), .b(net251) );
    and2_1 \U34_6_/U8  ( .x(\net225[9] ), .a(addr[6]), .b(net251) );
    and2_1 \U34_7_/U8  ( .x(\net225[8] ), .a(addr[7]), .b(net251) );
    and2_1 \U34_8_/U8  ( .x(\net225[7] ), .a(addr[32]), .b(net251) );
    and2_1 \U34_9_/U8  ( .x(\net225[6] ), .a(addr[33]), .b(net251) );
    and2_1 \U34_10_/U8  ( .x(\net225[5] ), .a(addr[34]), .b(net251) );
    and2_1 \U34_11_/U8  ( .x(\net225[4] ), .a(addr[35]), .b(net251) );
    and2_1 \U34_12_/U8  ( .x(\net225[3] ), .a(addr[36]), .b(net251) );
    and2_1 \U34_13_/U8  ( .x(\net225[2] ), .a(addr[37]), .b(net251) );
    and2_1 \U34_14_/U8  ( .x(\net225[1] ), .a(addr[38]), .b(net251) );
    and2_1 \U34_15_/U8  ( .x(\net225[0] ), .a(addr[39]), .b(net251) );
    and2_1 \U30_0_/U8  ( .x(\net222[15] ), .a(addr[24]), .b(net261) );
    and2_1 \U30_1_/U8  ( .x(\net222[14] ), .a(addr[25]), .b(net261) );
    and2_1 \U30_2_/U8  ( .x(\net222[13] ), .a(addr[26]), .b(net261) );
    and2_1 \U30_3_/U8  ( .x(\net222[12] ), .a(addr[27]), .b(net261) );
    and2_1 \U30_4_/U8  ( .x(\net222[11] ), .a(addr[28]), .b(net261) );
    and2_1 \U30_5_/U8  ( .x(\net222[10] ), .a(addr[29]), .b(net261) );
    and2_1 \U30_6_/U8  ( .x(\net222[9] ), .a(addr[30]), .b(net261) );
    and2_1 \U30_7_/U8  ( .x(\net222[8] ), .a(addr[31]), .b(net261) );
    and2_1 \U30_8_/U8  ( .x(\net222[7] ), .a(addr[56]), .b(net261) );
    and2_1 \U30_9_/U8  ( .x(\net222[6] ), .a(addr[57]), .b(net261) );
    and2_1 \U30_10_/U8  ( .x(\net222[5] ), .a(addr[58]), .b(net261) );
    and2_1 \U30_11_/U8  ( .x(\net222[4] ), .a(addr[59]), .b(net261) );
    and2_1 \U30_12_/U8  ( .x(\net222[3] ), .a(addr[60]), .b(net261) );
    and2_1 \U30_13_/U8  ( .x(\net222[2] ), .a(addr[61]), .b(net261) );
    and2_1 \U30_14_/U8  ( .x(\net222[1] ), .a(addr[62]), .b(net261) );
    and2_1 \U30_15_/U8  ( .x(\net222[0] ), .a(addr[63]), .b(net261) );
    and2_1 \U82_0_/U8  ( .x(\net219[15] ), .a(wd[0]), .b(net249) );
    and2_1 \U82_1_/U8  ( .x(\net219[14] ), .a(wd[1]), .b(net249) );
    and2_1 \U82_2_/U8  ( .x(\net219[13] ), .a(wd[2]), .b(net249) );
    and2_1 \U82_3_/U8  ( .x(\net219[12] ), .a(wd[3]), .b(net249) );
    and2_1 \U82_4_/U8  ( .x(\net219[11] ), .a(wd[4]), .b(net249) );
    and2_1 \U82_5_/U8  ( .x(\net219[10] ), .a(wd[5]), .b(net249) );
    and2_1 \U82_6_/U8  ( .x(\net219[9] ), .a(wd[6]), .b(net249) );
    and2_1 \U82_7_/U8  ( .x(\net219[8] ), .a(wd[7]), .b(net249) );
    and2_1 \U82_8_/U8  ( .x(\net219[7] ), .a(wd[32]), .b(net249) );
    and2_1 \U82_9_/U8  ( .x(\net219[6] ), .a(wd[33]), .b(net249) );
    and2_1 \U82_10_/U8  ( .x(\net219[5] ), .a(wd[34]), .b(net249) );
    and2_1 \U82_11_/U8  ( .x(\net219[4] ), .a(wd[35]), .b(net249) );
    and2_1 \U82_12_/U8  ( .x(\net219[3] ), .a(wd[36]), .b(net249) );
    and2_1 \U82_13_/U8  ( .x(\net219[2] ), .a(wd[37]), .b(net249) );
    and2_1 \U82_14_/U8  ( .x(\net219[1] ), .a(wd[38]), .b(net249) );
    and2_1 \U82_15_/U8  ( .x(\net219[0] ), .a(wd[39]), .b(net249) );
    inv_1 \U40_0_/U3  ( .x(\U40_0_/n3 ), .a(\net225[15] ) );
    inv_1 \U40_0_/U4  ( .x(\U40_0_/n4 ), .a(\net234[15] ) );
    inv_1 \U40_0_/U5  ( .x(\net217[15] ), .a(\U40_0_/n5 ) );
    inv_1 \U40_1_/U3  ( .x(\U40_1_/n3 ), .a(\net225[14] ) );
    inv_1 \U40_1_/U4  ( .x(\U40_1_/n4 ), .a(\net234[14] ) );
    inv_1 \U40_1_/U5  ( .x(\net217[14] ), .a(\U40_1_/n5 ) );
    inv_1 \U40_2_/U3  ( .x(\U40_2_/n3 ), .a(\net225[13] ) );
    inv_1 \U40_2_/U4  ( .x(\U40_2_/n4 ), .a(\net234[13] ) );
    inv_1 \U40_2_/U5  ( .x(\net217[13] ), .a(\U40_2_/n5 ) );
    inv_1 \U40_3_/U3  ( .x(\U40_3_/n3 ), .a(\net225[12] ) );
    inv_1 \U40_3_/U4  ( .x(\U40_3_/n4 ), .a(\net234[12] ) );
    inv_1 \U40_3_/U5  ( .x(\net217[12] ), .a(\U40_3_/n5 ) );
    inv_1 \U40_4_/U3  ( .x(\U40_4_/n3 ), .a(\net225[11] ) );
    inv_1 \U40_4_/U4  ( .x(\U40_4_/n4 ), .a(\net234[11] ) );
    inv_1 \U40_4_/U5  ( .x(\net217[11] ), .a(\U40_4_/n5 ) );
    inv_1 \U40_5_/U3  ( .x(\U40_5_/n3 ), .a(\net225[10] ) );
    inv_1 \U40_5_/U4  ( .x(\U40_5_/n4 ), .a(\net234[10] ) );
    inv_1 \U40_5_/U5  ( .x(\net217[10] ), .a(\U40_5_/n5 ) );
    inv_1 \U40_6_/U3  ( .x(\U40_6_/n3 ), .a(\net225[9] ) );
    inv_1 \U40_6_/U4  ( .x(\U40_6_/n4 ), .a(\net234[9] ) );
    inv_1 \U40_6_/U5  ( .x(\net217[9] ), .a(\U40_6_/n5 ) );
    inv_1 \U40_7_/U3  ( .x(\U40_7_/n3 ), .a(\net225[8] ) );
    inv_1 \U40_7_/U4  ( .x(\U40_7_/n4 ), .a(\net234[8] ) );
    inv_1 \U40_7_/U5  ( .x(\net217[8] ), .a(\U40_7_/n5 ) );
    inv_1 \U40_8_/U3  ( .x(\U40_8_/n3 ), .a(\net225[7] ) );
    inv_1 \U40_8_/U4  ( .x(\U40_8_/n4 ), .a(\net234[7] ) );
    inv_1 \U40_8_/U5  ( .x(\net217[7] ), .a(\U40_8_/n5 ) );
    inv_1 \U40_9_/U3  ( .x(\U40_9_/n3 ), .a(\net225[6] ) );
    inv_1 \U40_9_/U4  ( .x(\U40_9_/n4 ), .a(\net234[6] ) );
    inv_1 \U40_9_/U5  ( .x(\net217[6] ), .a(\U40_9_/n5 ) );
    inv_1 \U40_10_/U3  ( .x(\U40_10_/n3 ), .a(\net225[5] ) );
    inv_1 \U40_10_/U4  ( .x(\U40_10_/n4 ), .a(\net234[5] ) );
    inv_1 \U40_10_/U5  ( .x(\net217[5] ), .a(\U40_10_/n5 ) );
    inv_1 \U40_11_/U3  ( .x(\U40_11_/n3 ), .a(\net225[4] ) );
    inv_1 \U40_11_/U4  ( .x(\U40_11_/n4 ), .a(\net234[4] ) );
    inv_1 \U40_11_/U5  ( .x(\net217[4] ), .a(\U40_11_/n5 ) );
    inv_1 \U40_12_/U3  ( .x(\U40_12_/n3 ), .a(\net225[3] ) );
    inv_1 \U40_12_/U4  ( .x(\U40_12_/n4 ), .a(\net234[3] ) );
    inv_1 \U40_12_/U5  ( .x(\net217[3] ), .a(\U40_12_/n5 ) );
    inv_1 \U40_13_/U3  ( .x(\U40_13_/n3 ), .a(\net225[2] ) );
    inv_1 \U40_13_/U4  ( .x(\U40_13_/n4 ), .a(\net234[2] ) );
    inv_1 \U40_13_/U5  ( .x(\net217[2] ), .a(\U40_13_/n5 ) );
    inv_1 \U40_14_/U3  ( .x(\U40_14_/n3 ), .a(\net225[1] ) );
    inv_1 \U40_14_/U4  ( .x(\U40_14_/n4 ), .a(\net234[1] ) );
    inv_1 \U40_14_/U5  ( .x(\net217[1] ), .a(\U40_14_/n5 ) );
    inv_1 \U40_15_/U3  ( .x(\U40_15_/n3 ), .a(\net225[0] ) );
    inv_1 \U40_15_/U4  ( .x(\U40_15_/n4 ), .a(\net234[0] ) );
    inv_1 \U40_15_/U5  ( .x(\net217[0] ), .a(\U40_15_/n5 ) );
    and4_1 \U14_0_/U16  ( .x(\U14_0_/n5 ), .a(\U14_0_/n1 ), .b(\U14_0_/n2 ), 
        .c(\U14_0_/n3 ), .d(\U14_0_/n4 ) );
    inv_1 \U14_0_/U1  ( .x(\U14_0_/n1 ), .a(\net231[15] ) );
    inv_1 \U14_0_/U2  ( .x(\U14_0_/n2 ), .a(\net222[15] ) );
    inv_1 \U14_0_/U3  ( .x(\U14_0_/n3 ), .a(\net237[15] ) );
    inv_1 \U14_0_/U4  ( .x(\U14_0_/n4 ), .a(\net246[15] ) );
    inv_1 \U14_0_/U5  ( .x(\net212[15] ), .a(\U14_0_/n5 ) );
    and4_1 \U14_1_/U16  ( .x(\U14_1_/n5 ), .a(\U14_1_/n1 ), .b(\U14_1_/n2 ), 
        .c(\U14_1_/n3 ), .d(\U14_1_/n4 ) );
    inv_1 \U14_1_/U1  ( .x(\U14_1_/n1 ), .a(\net231[14] ) );
    inv_1 \U14_1_/U2  ( .x(\U14_1_/n2 ), .a(\net222[14] ) );
    inv_1 \U14_1_/U3  ( .x(\U14_1_/n3 ), .a(\net237[14] ) );
    inv_1 \U14_1_/U4  ( .x(\U14_1_/n4 ), .a(\net246[14] ) );
    inv_1 \U14_1_/U5  ( .x(\net212[14] ), .a(\U14_1_/n5 ) );
    and4_1 \U14_2_/U16  ( .x(\U14_2_/n5 ), .a(\U14_2_/n1 ), .b(\U14_2_/n2 ), 
        .c(\U14_2_/n3 ), .d(\U14_2_/n4 ) );
    inv_1 \U14_2_/U1  ( .x(\U14_2_/n1 ), .a(\net231[13] ) );
    inv_1 \U14_2_/U2  ( .x(\U14_2_/n2 ), .a(\net222[13] ) );
    inv_1 \U14_2_/U3  ( .x(\U14_2_/n3 ), .a(\net237[13] ) );
    inv_1 \U14_2_/U4  ( .x(\U14_2_/n4 ), .a(\net246[13] ) );
    inv_1 \U14_2_/U5  ( .x(\net212[13] ), .a(\U14_2_/n5 ) );
    and4_1 \U14_3_/U16  ( .x(\U14_3_/n5 ), .a(\U14_3_/n1 ), .b(\U14_3_/n2 ), 
        .c(\U14_3_/n3 ), .d(\U14_3_/n4 ) );
    inv_1 \U14_3_/U1  ( .x(\U14_3_/n1 ), .a(\net231[12] ) );
    inv_1 \U14_3_/U2  ( .x(\U14_3_/n2 ), .a(\net222[12] ) );
    inv_1 \U14_3_/U3  ( .x(\U14_3_/n3 ), .a(\net237[12] ) );
    inv_1 \U14_3_/U4  ( .x(\U14_3_/n4 ), .a(\net246[12] ) );
    inv_1 \U14_3_/U5  ( .x(\net212[12] ), .a(\U14_3_/n5 ) );
    and4_1 \U14_4_/U16  ( .x(\U14_4_/n5 ), .a(\U14_4_/n1 ), .b(\U14_4_/n2 ), 
        .c(\U14_4_/n3 ), .d(\U14_4_/n4 ) );
    inv_1 \U14_4_/U1  ( .x(\U14_4_/n1 ), .a(\net231[11] ) );
    inv_1 \U14_4_/U2  ( .x(\U14_4_/n2 ), .a(\net222[11] ) );
    inv_1 \U14_4_/U3  ( .x(\U14_4_/n3 ), .a(\net237[11] ) );
    inv_1 \U14_4_/U4  ( .x(\U14_4_/n4 ), .a(\net246[11] ) );
    inv_1 \U14_4_/U5  ( .x(\net212[11] ), .a(\U14_4_/n5 ) );
    and4_1 \U14_5_/U16  ( .x(\U14_5_/n5 ), .a(\U14_5_/n1 ), .b(\U14_5_/n2 ), 
        .c(\U14_5_/n3 ), .d(\U14_5_/n4 ) );
    inv_1 \U14_5_/U1  ( .x(\U14_5_/n1 ), .a(\net231[10] ) );
    inv_1 \U14_5_/U2  ( .x(\U14_5_/n2 ), .a(\net222[10] ) );
    inv_1 \U14_5_/U3  ( .x(\U14_5_/n3 ), .a(\net237[10] ) );
    inv_1 \U14_5_/U4  ( .x(\U14_5_/n4 ), .a(\net246[10] ) );
    inv_1 \U14_5_/U5  ( .x(\net212[10] ), .a(\U14_5_/n5 ) );
    and4_1 \U14_6_/U16  ( .x(\U14_6_/n5 ), .a(\U14_6_/n1 ), .b(\U14_6_/n2 ), 
        .c(\U14_6_/n3 ), .d(\U14_6_/n4 ) );
    inv_1 \U14_6_/U1  ( .x(\U14_6_/n1 ), .a(\net231[9] ) );
    inv_1 \U14_6_/U2  ( .x(\U14_6_/n2 ), .a(\net222[9] ) );
    inv_1 \U14_6_/U3  ( .x(\U14_6_/n3 ), .a(\net237[9] ) );
    inv_1 \U14_6_/U4  ( .x(\U14_6_/n4 ), .a(\net246[9] ) );
    inv_1 \U14_6_/U5  ( .x(\net212[9] ), .a(\U14_6_/n5 ) );
    and4_1 \U14_7_/U16  ( .x(\U14_7_/n5 ), .a(\U14_7_/n1 ), .b(\U14_7_/n2 ), 
        .c(\U14_7_/n3 ), .d(\U14_7_/n4 ) );
    inv_1 \U14_7_/U1  ( .x(\U14_7_/n1 ), .a(\net231[8] ) );
    inv_1 \U14_7_/U2  ( .x(\U14_7_/n2 ), .a(\net222[8] ) );
    inv_1 \U14_7_/U3  ( .x(\U14_7_/n3 ), .a(\net237[8] ) );
    inv_1 \U14_7_/U4  ( .x(\U14_7_/n4 ), .a(\net246[8] ) );
    inv_1 \U14_7_/U5  ( .x(\net212[8] ), .a(\U14_7_/n5 ) );
    and4_1 \U14_8_/U16  ( .x(\U14_8_/n5 ), .a(\U14_8_/n1 ), .b(\U14_8_/n2 ), 
        .c(\U14_8_/n3 ), .d(\U14_8_/n4 ) );
    inv_1 \U14_8_/U1  ( .x(\U14_8_/n1 ), .a(\net231[7] ) );
    inv_1 \U14_8_/U2  ( .x(\U14_8_/n2 ), .a(\net222[7] ) );
    inv_1 \U14_8_/U3  ( .x(\U14_8_/n3 ), .a(\net237[7] ) );
    inv_1 \U14_8_/U4  ( .x(\U14_8_/n4 ), .a(\net246[7] ) );
    inv_1 \U14_8_/U5  ( .x(\net212[7] ), .a(\U14_8_/n5 ) );
    and4_1 \U14_9_/U16  ( .x(\U14_9_/n5 ), .a(\U14_9_/n1 ), .b(\U14_9_/n2 ), 
        .c(\U14_9_/n3 ), .d(\U14_9_/n4 ) );
    inv_1 \U14_9_/U1  ( .x(\U14_9_/n1 ), .a(\net231[6] ) );
    inv_1 \U14_9_/U2  ( .x(\U14_9_/n2 ), .a(\net222[6] ) );
    inv_1 \U14_9_/U3  ( .x(\U14_9_/n3 ), .a(\net237[6] ) );
    inv_1 \U14_9_/U4  ( .x(\U14_9_/n4 ), .a(\net246[6] ) );
    inv_1 \U14_9_/U5  ( .x(\net212[6] ), .a(\U14_9_/n5 ) );
    and4_1 \U14_10_/U16  ( .x(\U14_10_/n5 ), .a(\U14_10_/n1 ), .b(\U14_10_/n2 
        ), .c(\U14_10_/n3 ), .d(\U14_10_/n4 ) );
    inv_1 \U14_10_/U1  ( .x(\U14_10_/n1 ), .a(\net231[5] ) );
    inv_1 \U14_10_/U2  ( .x(\U14_10_/n2 ), .a(\net222[5] ) );
    inv_1 \U14_10_/U3  ( .x(\U14_10_/n3 ), .a(\net237[5] ) );
    inv_1 \U14_10_/U4  ( .x(\U14_10_/n4 ), .a(\net246[5] ) );
    inv_1 \U14_10_/U5  ( .x(\net212[5] ), .a(\U14_10_/n5 ) );
    inv_1 \U14_11_/U1  ( .x(\U14_11_/n1 ), .a(\net231[4] ) );
    inv_1 \U14_11_/U2  ( .x(\U14_11_/n2 ), .a(\net222[4] ) );
    inv_1 \U14_11_/U4  ( .x(\U14_11_/n4 ), .a(\net246[4] ) );
    inv_1 \U14_11_/U5  ( .x(\net212[4] ), .a(\U14_11_/n5 ) );
    inv_1 \U14_12_/U1  ( .x(\U14_12_/n1 ), .a(\net231[3] ) );
    inv_1 \U14_12_/U2  ( .x(\U14_12_/n2 ), .a(\net222[3] ) );
    inv_1 \U14_12_/U4  ( .x(\U14_12_/n4 ), .a(\net246[3] ) );
    inv_1 \U14_12_/U5  ( .x(\net212[3] ), .a(\U14_12_/n5 ) );
    and4_1 \U14_13_/U16  ( .x(\U14_13_/n5 ), .a(\U14_13_/n1 ), .b(\U14_13_/n2 
        ), .c(\U14_13_/n3 ), .d(\U14_13_/n4 ) );
    inv_1 \U14_13_/U1  ( .x(\U14_13_/n1 ), .a(\net231[2] ) );
    inv_1 \U14_13_/U2  ( .x(\U14_13_/n2 ), .a(\net222[2] ) );
    inv_1 \U14_13_/U3  ( .x(\U14_13_/n3 ), .a(\net237[2] ) );
    inv_1 \U14_13_/U4  ( .x(\U14_13_/n4 ), .a(\net246[2] ) );
    inv_1 \U14_13_/U5  ( .x(\net212[2] ), .a(\U14_13_/n5 ) );
    and4_1 \U14_14_/U16  ( .x(\U14_14_/n5 ), .a(\U14_14_/n1 ), .b(\U14_14_/n2 
        ), .c(\U14_14_/n3 ), .d(\U14_14_/n4 ) );
    inv_1 \U14_14_/U1  ( .x(\U14_14_/n1 ), .a(\net231[1] ) );
    inv_1 \U14_14_/U2  ( .x(\U14_14_/n2 ), .a(\net222[1] ) );
    inv_1 \U14_14_/U3  ( .x(\U14_14_/n3 ), .a(\net237[1] ) );
    inv_1 \U14_14_/U4  ( .x(\U14_14_/n4 ), .a(\net246[1] ) );
    inv_1 \U14_14_/U5  ( .x(\net212[1] ), .a(\U14_14_/n5 ) );
    and4_1 \U14_15_/U16  ( .x(\U14_15_/n5 ), .a(\U14_15_/n1 ), .b(\U14_15_/n2 
        ), .c(\U14_15_/n3 ), .d(\U14_15_/n4 ) );
    inv_1 \U14_15_/U1  ( .x(\U14_15_/n1 ), .a(\net231[0] ) );
    inv_1 \U14_15_/U2  ( .x(\U14_15_/n2 ), .a(\net222[0] ) );
    inv_1 \U14_15_/U3  ( .x(\U14_15_/n3 ), .a(\net237[0] ) );
    inv_1 \U14_15_/U4  ( .x(\U14_15_/n4 ), .a(\net246[0] ) );
    inv_1 \U14_15_/U5  ( .x(\net212[0] ), .a(\U14_15_/n5 ) );
    and4_1 \U91_0_/U16  ( .x(\U91_0_/n5 ), .a(\U91_0_/n1 ), .b(\U91_0_/n2 ), 
        .c(\U91_0_/n3 ), .d(\U91_0_/n4 ) );
    inv_1 \U91_0_/U1  ( .x(\U91_0_/n1 ), .a(\net219[15] ) );
    inv_1 \U91_0_/U2  ( .x(\U91_0_/n2 ), .a(\net243[15] ) );
    inv_1 \U91_0_/U3  ( .x(\U91_0_/n3 ), .a(\net240[15] ) );
    inv_1 \U91_0_/U4  ( .x(\U91_0_/n4 ), .a(\net228[15] ) );
    inv_1 \U91_0_/U5  ( .x(\net207[15] ), .a(\U91_0_/n5 ) );
    and4_1 \U91_1_/U16  ( .x(\U91_1_/n5 ), .a(\U91_1_/n1 ), .b(\U91_1_/n2 ), 
        .c(\U91_1_/n3 ), .d(\U91_1_/n4 ) );
    inv_1 \U91_1_/U1  ( .x(\U91_1_/n1 ), .a(\net219[14] ) );
    inv_1 \U91_1_/U2  ( .x(\U91_1_/n2 ), .a(\net243[14] ) );
    inv_1 \U91_1_/U3  ( .x(\U91_1_/n3 ), .a(\net240[14] ) );
    inv_1 \U91_1_/U4  ( .x(\U91_1_/n4 ), .a(\net228[14] ) );
    inv_1 \U91_1_/U5  ( .x(\net207[14] ), .a(\U91_1_/n5 ) );
    and4_1 \U91_2_/U16  ( .x(\U91_2_/n5 ), .a(\U91_2_/n1 ), .b(\U91_2_/n2 ), 
        .c(\U91_2_/n3 ), .d(\U91_2_/n4 ) );
    inv_1 \U91_2_/U1  ( .x(\U91_2_/n1 ), .a(\net219[13] ) );
    inv_1 \U91_2_/U2  ( .x(\U91_2_/n2 ), .a(\net243[13] ) );
    inv_1 \U91_2_/U3  ( .x(\U91_2_/n3 ), .a(\net240[13] ) );
    inv_1 \U91_2_/U4  ( .x(\U91_2_/n4 ), .a(\net228[13] ) );
    inv_1 \U91_2_/U5  ( .x(\net207[13] ), .a(\U91_2_/n5 ) );
    and4_1 \U91_3_/U16  ( .x(\U91_3_/n5 ), .a(\U91_3_/n1 ), .b(\U91_3_/n2 ), 
        .c(\U91_3_/n3 ), .d(\U91_3_/n4 ) );
    inv_1 \U91_3_/U1  ( .x(\U91_3_/n1 ), .a(\net219[12] ) );
    inv_1 \U91_3_/U2  ( .x(\U91_3_/n2 ), .a(\net243[12] ) );
    inv_1 \U91_3_/U3  ( .x(\U91_3_/n3 ), .a(\net240[12] ) );
    inv_1 \U91_3_/U4  ( .x(\U91_3_/n4 ), .a(\net228[12] ) );
    inv_1 \U91_3_/U5  ( .x(\net207[12] ), .a(\U91_3_/n5 ) );
    and4_1 \U91_4_/U16  ( .x(\U91_4_/n5 ), .a(\U91_4_/n1 ), .b(\U91_4_/n2 ), 
        .c(\U91_4_/n3 ), .d(\U91_4_/n4 ) );
    inv_1 \U91_4_/U1  ( .x(\U91_4_/n1 ), .a(\net219[11] ) );
    inv_1 \U91_4_/U2  ( .x(\U91_4_/n2 ), .a(\net243[11] ) );
    inv_1 \U91_4_/U3  ( .x(\U91_4_/n3 ), .a(\net240[11] ) );
    inv_1 \U91_4_/U4  ( .x(\U91_4_/n4 ), .a(\net228[11] ) );
    inv_1 \U91_4_/U5  ( .x(\net207[11] ), .a(\U91_4_/n5 ) );
    and4_1 \U91_5_/U16  ( .x(\U91_5_/n5 ), .a(\U91_5_/n1 ), .b(\U91_5_/n2 ), 
        .c(\U91_5_/n3 ), .d(\U91_5_/n4 ) );
    inv_1 \U91_5_/U1  ( .x(\U91_5_/n1 ), .a(\net219[10] ) );
    inv_1 \U91_5_/U2  ( .x(\U91_5_/n2 ), .a(\net243[10] ) );
    inv_1 \U91_5_/U3  ( .x(\U91_5_/n3 ), .a(\net240[10] ) );
    inv_1 \U91_5_/U4  ( .x(\U91_5_/n4 ), .a(\net228[10] ) );
    inv_1 \U91_5_/U5  ( .x(\net207[10] ), .a(\U91_5_/n5 ) );
    and4_1 \U91_6_/U16  ( .x(\U91_6_/n5 ), .a(\U91_6_/n1 ), .b(\U91_6_/n2 ), 
        .c(\U91_6_/n3 ), .d(\U91_6_/n4 ) );
    inv_1 \U91_6_/U1  ( .x(\U91_6_/n1 ), .a(\net219[9] ) );
    inv_1 \U91_6_/U2  ( .x(\U91_6_/n2 ), .a(\net243[9] ) );
    inv_1 \U91_6_/U3  ( .x(\U91_6_/n3 ), .a(\net240[9] ) );
    inv_1 \U91_6_/U4  ( .x(\U91_6_/n4 ), .a(\net228[9] ) );
    inv_1 \U91_6_/U5  ( .x(\net207[9] ), .a(\U91_6_/n5 ) );
    and4_1 \U91_7_/U16  ( .x(\U91_7_/n5 ), .a(\U91_7_/n1 ), .b(\U91_7_/n2 ), 
        .c(\U91_7_/n3 ), .d(\U91_7_/n4 ) );
    inv_1 \U91_7_/U1  ( .x(\U91_7_/n1 ), .a(\net219[8] ) );
    inv_1 \U91_7_/U2  ( .x(\U91_7_/n2 ), .a(\net243[8] ) );
    inv_1 \U91_7_/U3  ( .x(\U91_7_/n3 ), .a(\net240[8] ) );
    inv_1 \U91_7_/U4  ( .x(\U91_7_/n4 ), .a(\net228[8] ) );
    inv_1 \U91_7_/U5  ( .x(\net207[8] ), .a(\U91_7_/n5 ) );
    and4_1 \U91_8_/U16  ( .x(\U91_8_/n5 ), .a(\U91_8_/n1 ), .b(\U91_8_/n2 ), 
        .c(\U91_8_/n3 ), .d(\U91_8_/n4 ) );
    inv_1 \U91_8_/U1  ( .x(\U91_8_/n1 ), .a(\net219[7] ) );
    inv_1 \U91_8_/U2  ( .x(\U91_8_/n2 ), .a(\net243[7] ) );
    inv_1 \U91_8_/U3  ( .x(\U91_8_/n3 ), .a(\net240[7] ) );
    inv_1 \U91_8_/U4  ( .x(\U91_8_/n4 ), .a(\net228[7] ) );
    inv_1 \U91_8_/U5  ( .x(\net207[7] ), .a(\U91_8_/n5 ) );
    and4_1 \U91_9_/U16  ( .x(\U91_9_/n5 ), .a(\U91_9_/n1 ), .b(\U91_9_/n2 ), 
        .c(\U91_9_/n3 ), .d(\U91_9_/n4 ) );
    inv_1 \U91_9_/U1  ( .x(\U91_9_/n1 ), .a(\net219[6] ) );
    inv_1 \U91_9_/U2  ( .x(\U91_9_/n2 ), .a(\net243[6] ) );
    inv_1 \U91_9_/U3  ( .x(\U91_9_/n3 ), .a(\net240[6] ) );
    inv_1 \U91_9_/U4  ( .x(\U91_9_/n4 ), .a(\net228[6] ) );
    inv_1 \U91_9_/U5  ( .x(\net207[6] ), .a(\U91_9_/n5 ) );
    and4_1 \U91_10_/U16  ( .x(\U91_10_/n5 ), .a(\U91_10_/n1 ), .b(\U91_10_/n2 
        ), .c(\U91_10_/n3 ), .d(\U91_10_/n4 ) );
    inv_1 \U91_10_/U1  ( .x(\U91_10_/n1 ), .a(\net219[5] ) );
    inv_1 \U91_10_/U2  ( .x(\U91_10_/n2 ), .a(\net243[5] ) );
    inv_1 \U91_10_/U3  ( .x(\U91_10_/n3 ), .a(\net240[5] ) );
    inv_1 \U91_10_/U4  ( .x(\U91_10_/n4 ), .a(\net228[5] ) );
    inv_1 \U91_10_/U5  ( .x(\net207[5] ), .a(\U91_10_/n5 ) );
    and4_1 \U91_11_/U16  ( .x(\U91_11_/n5 ), .a(\U91_11_/n1 ), .b(\U91_11_/n2 
        ), .c(\U91_11_/n3 ), .d(\U91_11_/n4 ) );
    inv_1 \U91_11_/U1  ( .x(\U91_11_/n1 ), .a(\net219[4] ) );
    inv_1 \U91_11_/U2  ( .x(\U91_11_/n2 ), .a(\net243[4] ) );
    inv_1 \U91_11_/U3  ( .x(\U91_11_/n3 ), .a(\net240[4] ) );
    inv_1 \U91_11_/U4  ( .x(\U91_11_/n4 ), .a(\net228[4] ) );
    inv_1 \U91_11_/U5  ( .x(\net207[4] ), .a(\U91_11_/n5 ) );
    and4_1 \U91_12_/U16  ( .x(\U91_12_/n5 ), .a(\U91_12_/n1 ), .b(\U91_12_/n2 
        ), .c(\U91_12_/n3 ), .d(\U91_12_/n4 ) );
    inv_1 \U91_12_/U1  ( .x(\U91_12_/n1 ), .a(\net219[3] ) );
    inv_1 \U91_12_/U2  ( .x(\U91_12_/n2 ), .a(\net243[3] ) );
    inv_1 \U91_12_/U3  ( .x(\U91_12_/n3 ), .a(\net240[3] ) );
    inv_1 \U91_12_/U4  ( .x(\U91_12_/n4 ), .a(\net228[3] ) );
    inv_1 \U91_12_/U5  ( .x(\net207[3] ), .a(\U91_12_/n5 ) );
    and4_1 \U91_13_/U16  ( .x(\U91_13_/n5 ), .a(\U91_13_/n1 ), .b(\U91_13_/n2 
        ), .c(\U91_13_/n3 ), .d(\U91_13_/n4 ) );
    inv_1 \U91_13_/U1  ( .x(\U91_13_/n1 ), .a(\net219[2] ) );
    inv_1 \U91_13_/U2  ( .x(\U91_13_/n2 ), .a(\net243[2] ) );
    inv_1 \U91_13_/U3  ( .x(\U91_13_/n3 ), .a(\net240[2] ) );
    inv_1 \U91_13_/U4  ( .x(\U91_13_/n4 ), .a(\net228[2] ) );
    inv_1 \U91_13_/U5  ( .x(\net207[2] ), .a(\U91_13_/n5 ) );
    and4_1 \U91_14_/U16  ( .x(\U91_14_/n5 ), .a(\U91_14_/n1 ), .b(\U91_14_/n2 
        ), .c(\U91_14_/n3 ), .d(\U91_14_/n4 ) );
    inv_1 \U91_14_/U1  ( .x(\U91_14_/n1 ), .a(\net219[1] ) );
    inv_1 \U91_14_/U2  ( .x(\U91_14_/n2 ), .a(\net243[1] ) );
    inv_1 \U91_14_/U3  ( .x(\U91_14_/n3 ), .a(\net240[1] ) );
    inv_1 \U91_14_/U4  ( .x(\U91_14_/n4 ), .a(\net228[1] ) );
    inv_1 \U91_14_/U5  ( .x(\net207[1] ), .a(\U91_14_/n5 ) );
    and4_1 \U91_15_/U16  ( .x(\U91_15_/n5 ), .a(\U91_15_/n1 ), .b(\U91_15_/n2 
        ), .c(\U91_15_/n3 ), .d(\U91_15_/n4 ) );
    inv_1 \U91_15_/U1  ( .x(\U91_15_/n1 ), .a(\net219[0] ) );
    inv_1 \U91_15_/U2  ( .x(\U91_15_/n2 ), .a(\net243[0] ) );
    inv_1 \U91_15_/U3  ( .x(\U91_15_/n3 ), .a(\net240[0] ) );
    inv_1 \U91_15_/U4  ( .x(\U91_15_/n4 ), .a(\net228[0] ) );
    inv_1 \U91_15_/U5  ( .x(\net207[0] ), .a(\U91_15_/n5 ) );
    or3_2 \U93_0_/U12  ( .x(chainl[0]), .a(\net207[15] ), .b(\net217[15] ), 
        .c(\net212[15] ) );
    or3_2 \U93_1_/U12  ( .x(chainl[1]), .a(\net207[14] ), .b(\net217[14] ), 
        .c(\net212[14] ) );
    or3_2 \U93_2_/U12  ( .x(chainl[2]), .a(\net207[13] ), .b(\net217[13] ), 
        .c(\net212[13] ) );
    or3_2 \U93_3_/U12  ( .x(chainl[3]), .a(\net207[12] ), .b(\net217[12] ), 
        .c(\net212[12] ) );
    or3_2 \U93_4_/U12  ( .x(chainl[4]), .a(\net207[11] ), .b(\net217[11] ), 
        .c(\net212[11] ) );
    or3_2 \U93_5_/U12  ( .x(chainl[5]), .a(\net207[10] ), .b(\net217[10] ), 
        .c(\net212[10] ) );
    or3_2 \U93_6_/U12  ( .x(chainl[6]), .a(\net207[9] ), .b(\net217[9] ), .c(
        \net212[9] ) );
    or3_2 \U93_7_/U12  ( .x(chainl[7]), .a(\net207[8] ), .b(\net217[8] ), .c(
        \net212[8] ) );
    or3_2 \U93_8_/U12  ( .x(chainh[0]), .a(\net207[7] ), .b(\net217[7] ), .c(
        \net212[7] ) );
    or3_2 \U93_9_/U12  ( .x(chainh[1]), .a(\net207[6] ), .b(\net217[6] ), .c(
        \net212[6] ) );
    or3_2 \U93_10_/U12  ( .x(chainh[2]), .a(\net207[5] ), .b(\net217[5] ), .c(
        \net212[5] ) );
    or3_2 \U93_11_/U12  ( .x(chainh[3]), .a(\net207[4] ), .b(\net217[4] ), .c(
        \net212[4] ) );
    or3_2 \U93_12_/U12  ( .x(chainh[4]), .a(\net207[3] ), .b(\net217[3] ), .c(
        \net212[3] ) );
    or3_2 \U93_13_/U12  ( .x(chainh[5]), .a(\net207[2] ), .b(\net217[2] ), .c(
        \net212[2] ) );
    or3_2 \U93_14_/U12  ( .x(chainh[6]), .a(\net207[1] ), .b(\net217[1] ), .c(
        \net212[1] ) );
    or3_2 \U93_15_/U12  ( .x(chainh[7]), .a(\net207[0] ), .b(\net217[0] ), .c(
        \net212[0] ) );
    inv_1 \U152/U3  ( .x(net198), .a(sendreq) );
    ao23_1 \U158/U19/U21/U1/U1  ( .x(net131), .a(net132), .b(net131), .c(
        net132), .d(rnw[1]), .e(rnw[1]) );
    ao23_1 \U157/U19/U21/U1/U1  ( .x(net176), .a(net132), .b(net176), .c(
        net132), .d(rnw[0]), .e(rnw[0]) );
    ao222_1 \U123/U18/U1/U1  ( .x(net136), .a(net185), .b(net187), .c(net185), 
        .d(net136), .e(net187), .f(net136) );
    aoi21_1 \U151/U30/U1/U1  ( .x(\hdr[4] ), .a(\U151/Z ), .b(net138), .c(
        net198) );
    inv_1 \U151/U30/U1/U2  ( .x(\U151/Z ), .a(\hdr[4] ) );
    nor3_1 \U148/U21/Unr  ( .x(\U148/U21/nr ), .a(net191), .b(net136), .c(
        net293) );
    nand3_1 \U148/U21/Und  ( .x(\U148/U21/nd ), .a(net191), .b(net136), .c(
        net293) );
    oa21_1 \U148/U21/U1  ( .x(\U148/U21/n2 ), .a(\U148/U21/n2 ), .b(
        \U148/U21/nr ), .c(\U148/U21/nd ) );
    inv_1 \U148/U21/U3  ( .x(ack), .a(\U148/U21/n2 ) );
    buf_3 U1 ( .x(n1), .a(net138) );
    buf_3 U2 ( .x(net138), .a(nia) );
    buf_3 U3 ( .x(net269), .a(net146) );
    buf_3 U4 ( .x(net255), .a(\bs[5] ) );
    buf_3 U5 ( .x(net267), .a(\bs[6] ) );
    buf_3 U6 ( .x(net263), .a(\bs[7] ) );
    buf_3 U7 ( .x(net249), .a(\bs[8] ) );
    buf_3 U8 ( .x(net253), .a(\bs[2] ) );
    buf_3 U9 ( .x(net251), .a(\bs[4] ) );
    buf_3 U10 ( .x(net259), .a(\bs[3] ) );
    buf_3 U11 ( .x(net261), .a(\bs[1] ) );
    buf_3 U12 ( .x(net265), .a(\bs[0] ) );
    and2_1 U13 ( .x(\U40_2_/n5 ), .a(\U40_2_/n3 ), .b(\U40_2_/n4 ) );
    and2_1 U14 ( .x(\U40_1_/n5 ), .a(\U40_1_/n3 ), .b(\U40_1_/n4 ) );
    and2_1 U15 ( .x(\U40_9_/n5 ), .a(\U40_9_/n3 ), .b(\U40_9_/n4 ) );
    and2_1 U16 ( .x(\U40_8_/n5 ), .a(\U40_8_/n3 ), .b(\U40_8_/n4 ) );
    and2_1 U17 ( .x(\U40_13_/n5 ), .a(\U40_13_/n3 ), .b(\U40_13_/n4 ) );
    and2_1 U18 ( .x(\U40_0_/n5 ), .a(\U40_0_/n3 ), .b(\U40_0_/n4 ) );
    and2_1 U19 ( .x(\U40_5_/n5 ), .a(\U40_5_/n3 ), .b(\U40_5_/n4 ) );
    and2_1 U20 ( .x(\U40_4_/n5 ), .a(\U40_4_/n3 ), .b(\U40_4_/n4 ) );
    and3_1 U21 ( .x(\U14_12_/n5 ), .a(\U14_12_/n2 ), .b(\U14_12_/n4 ), .c(
        \U14_12_/n1 ) );
    and2_1 U22 ( .x(\U40_12_/n5 ), .a(\U40_12_/n3 ), .b(\U40_12_/n4 ) );
    and2_1 U23 ( .x(\U40_3_/n5 ), .a(\U40_3_/n3 ), .b(\U40_3_/n4 ) );
    and3_1 U24 ( .x(\U14_11_/n5 ), .a(\U14_11_/n2 ), .b(\U14_11_/n4 ), .c(
        \U14_11_/n1 ) );
    and2_1 U25 ( .x(\U40_11_/n5 ), .a(\U40_11_/n3 ), .b(\U40_11_/n4 ) );
    and2_1 U26 ( .x(\U40_10_/n5 ), .a(\U40_10_/n3 ), .b(\U40_10_/n4 ) );
    and2_1 U27 ( .x(\U40_15_/n5 ), .a(\U40_15_/n3 ), .b(\U40_15_/n4 ) );
    and2_1 U28 ( .x(\U40_7_/n5 ), .a(\U40_7_/n3 ), .b(\U40_7_/n4 ) );
    and2_1 U29 ( .x(\U40_6_/n5 ), .a(\U40_6_/n3 ), .b(\U40_6_/n4 ) );
    and2_1 U30 ( .x(\U40_14_/n5 ), .a(\U40_14_/n3 ), .b(\U40_14_/n4 ) );
endmodule


module chain_ic_ctrl_1 ( ack, candefer, eop, nstatack, pltxreq, routetxreq, 
    tok_ack, accept, candefer_ack, defer, eopack, lock, nReset, pltxack, 
    routetxack, tok_err, tok_ok );
input  [1:0] candefer_ack;
input  [1:0] lock;
input  accept, defer, eopack, nReset, pltxack, routetxack, tok_err, tok_ok;
output ack, candefer, eop, nstatack, pltxreq, routetxreq, tok_ack;
    wire \locked[1] , \locked[0] , net21, net12, net20, net16, net10, net7, 
        net6, retry, net27, txnodefer, net13, txunlocked, net5, txmaydefer, 
        txdone, net8, txlocked, net29, net2, net4, lockcleared, net28, net18, 
        net22, net14, net9, net24, net19, net31, net11, net30, net17, net3, 
        reset, net26, nlclear, lwrite, net15, net23, net25, \U249/n5 , 
        \U249/n1 , \U249/n2 , \U249/n3 , \U249/n4 , \U286/U28/U1/clr , 
        \U286/U28/U1/set , \U285/U28/U1/clr , \U285/U28/U1/set , 
        \U262/U25/U1/clr , \U262/U25/U1/ob , \U284/U25/U1/clr , 
        \U284/U25/U1/ob , \U283/U25/U1/clr , \U283/U25/U1/ob , \U288/Z , 
        \U289/Z , \U287/Z , \U149/nr , \U149/nd , \U149/n2 , \U160/acb , 
        \U160/U1/Z , \U136/nlsense , \U136/nulsense , \U136/nwh , \U136/nwl , 
        \U136/nclear_latch , n1, n2;
    nand2_1 \U146/U5  ( .x(candefer), .a(net23), .b(net25) );
    or2_1 \U277/U12  ( .x(net6), .a(net19), .b(net9) );
    or2_1 \U264/U12  ( .x(retry), .a(net31), .b(net24) );
    or2_1 \U259/U12  ( .x(net28), .a(net27), .b(net7) );
    or2_1 \U140/U12  ( .x(net18), .a(net13), .b(net8) );
    or2_1 \U148/U12  ( .x(net11), .a(net15), .b(routetxack) );
    and4_1 \U249/U16  ( .x(\U249/n5 ), .a(\U249/n1 ), .b(\U249/n2 ), .c(
        \U249/n3 ), .d(\U249/n4 ) );
    inv_1 \U249/U1  ( .x(\U249/n1 ), .a(txnodefer) );
    inv_1 \U249/U2  ( .x(\U249/n2 ), .a(net16) );
    inv_1 \U249/U3  ( .x(\U249/n3 ), .a(net9) );
    inv_1 \U249/U4  ( .x(\U249/n4 ), .a(net19) );
    inv_1 \U249/U5  ( .x(ack), .a(\U249/n5 ) );
    nor3_2 \U40/U16  ( .x(nstatack), .a(net16), .b(reset), .c(retry) );
    nor3_2 \U275/U16  ( .x(net17), .a(net29), .b(reset), .c(tok_ack) );
    buf_3 \U290/U8  ( .x(net12), .a(txmaydefer) );
    nor2_1 \U154/U5  ( .x(nlclear), .a(net4), .b(net31) );
    or2_2 \U274/U12  ( .x(pltxreq), .a(net22), .b(net14) );
    or3_1 \U260/U12  ( .x(eop), .a(net31), .b(txlocked), .c(net4) );
    inv_1 \U147/U3  ( .x(net3), .a(net29) );
    inv_1 \U174/U3  ( .x(reset), .a(nReset) );
    aoai211_1 \U286/U28/U1/U1  ( .x(\U286/U28/U1/clr ), .a(net3), .b(n1), .c(
        net17), .d(net22) );
    nand3_1 \U286/U28/U1/U2  ( .x(\U286/U28/U1/set ), .a(net17), .b(net3), .c(
        n1) );
    nand2_2 \U286/U28/U1/U3  ( .x(net22), .a(\U286/U28/U1/clr ), .b(
        \U286/U28/U1/set ) );
    aoai211_1 \U285/U28/U1/U1  ( .x(\U285/U28/U1/clr ), .a(net3), .b(n2), .c(
        net17), .d(net14) );
    nand3_1 \U285/U28/U1/U2  ( .x(\U285/U28/U1/set ), .a(net17), .b(net3), .c(
        n2) );
    nand2_2 \U285/U28/U1/U3  ( .x(net14), .a(\U285/U28/U1/clr ), .b(
        \U285/U28/U1/set ) );
    ao222_1 \U254/U18/U1/U1  ( .x(net31), .a(defer), .b(txunlocked), .c(defer), 
        .d(net31), .e(txunlocked), .f(net31) );
    ao222_1 \U252/U18/U1/U1  ( .x(net19), .a(tok_err), .b(net12), .c(tok_err), 
        .d(net19), .e(net12), .f(net19) );
    ao222_1 \U276/U18/U1/U1  ( .x(net24), .a(txlocked), .b(defer), .c(txlocked
        ), .d(net24), .e(defer), .f(net24) );
    ao222_1 \U251/U18/U1/U1  ( .x(net9), .a(tok_ok), .b(net12), .c(tok_ok), 
        .d(net9), .e(net12), .f(net9) );
    ao222_1 \U235/U18/U1/U1  ( .x(tok_ack), .a(ack), .b(net2), .c(ack), .d(
        tok_ack), .e(net2), .f(tok_ack) );
    ao222_1 \U247/U18/U1/U1  ( .x(txnodefer), .a(txdone), .b(candefer_ack[0]), 
        .c(txdone), .d(txnodefer), .e(candefer_ack[0]), .f(txnodefer) );
    ao222_2 \U246/U19/U1/U1  ( .x(txlocked), .a(net14), .b(txdone), .c(net14), 
        .d(txlocked), .e(txdone), .f(txlocked) );
    ao222_2 \U245/U19/U1/U1  ( .x(txunlocked), .a(txdone), .b(net22), .c(
        txdone), .d(txunlocked), .e(net22), .f(txunlocked) );
    ao222_1 \U269/U18/U1/U1  ( .x(net2), .a(net28), .b(net18), .c(net28), .d(
        net2), .e(net18), .f(net2) );
    ao222_1 \U268/U18/U1/U1  ( .x(net5), .a(eopack), .b(lockcleared), .c(
        eopack), .d(net5), .e(lockcleared), .f(net5) );
    ao222_1 \U256/U18/U1/U1  ( .x(net4), .a(tok_err), .b(txunlocked), .c(
        tok_err), .d(net4), .e(txunlocked), .f(net4) );
    ao222_1 \U175/U18/U1/U1  ( .x(net29), .a(net2), .b(retry), .c(net2), .d(
        net29), .e(retry), .f(net29) );
    ao222_1 \U255/U18/U1/U1  ( .x(net8), .a(txlocked), .b(eopack), .c(txlocked
        ), .d(net8), .e(eopack), .f(net8) );
    ao222_2 \U248/U19/U1/U1  ( .x(txmaydefer), .a(candefer_ack[1]), .b(txdone), 
        .c(candefer_ack[1]), .d(txmaydefer), .e(txdone), .f(txmaydefer) );
    ao222_2 \U250/U19/U1/U1  ( .x(net16), .a(accept), .b(net12), .c(accept), 
        .d(net16), .e(net12), .f(net16) );
    oa31_1 \U262/U25/U1/Uclr  ( .x(\U262/U25/U1/clr ), .a(txunlocked), .b(net5
        ), .c(tok_ok), .d(net13) );
    oaoi211_1 \U262/U25/U1/Uaoi  ( .x(\U262/U25/U1/ob ), .a(net5), .b(tok_ok), 
        .c(txunlocked), .d(\U262/U25/U1/clr ) );
    inv_2 \U262/U25/U1/Ui  ( .x(net13), .a(\U262/U25/U1/ob ) );
    oa31_1 \U284/U25/U1/Uclr  ( .x(\U284/U25/U1/clr ), .a(txnodefer), .b(
        tok_ok), .c(tok_err), .d(net27) );
    oaoi211_1 \U284/U25/U1/Uaoi  ( .x(\U284/U25/U1/ob ), .a(tok_ok), .b(
        tok_err), .c(txnodefer), .d(\U284/U25/U1/clr ) );
    inv_2 \U284/U25/U1/Ui  ( .x(net27), .a(\U284/U25/U1/ob ) );
    oa31_1 \U283/U25/U1/Uclr  ( .x(\U283/U25/U1/clr ), .a(net10), .b(net6), 
        .c(retry), .d(net7) );
    oaoi211_1 \U283/U25/U1/Uaoi  ( .x(\U283/U25/U1/ob ), .a(net6), .b(retry), 
        .c(net10), .d(\U283/U25/U1/clr ) );
    inv_2 \U283/U25/U1/Ui  ( .x(net7), .a(\U283/U25/U1/ob ) );
    aoi21_1 \U289/U30/U1/U1  ( .x(net20), .a(\U289/Z ), .b(net16), .c(net12)
         );
    inv_1 \U289/U30/U1/U2  ( .x(\U289/Z ), .a(net20) );
    aoi21_1 \U287/U30/U1/U1  ( .x(net21), .a(\U287/Z ), .b(accept), .c(net12)
         );
    inv_1 \U287/U30/U1/U2  ( .x(\U287/Z ), .a(net21) );
    aoi222_1 \U288/U30/U1  ( .x(net10), .a(net20), .b(net21), .c(net20), .d(
        \U288/Z ), .e(net21), .f(\U288/Z ) );
    inv_1 \U288/U30/Uinv  ( .x(\U288/Z ), .a(net10) );
    nor3_1 \U149/Unr  ( .x(\U149/nr ), .a(pltxack), .b(net11), .c(net30) );
    nand3_1 \U149/Und  ( .x(\U149/nd ), .a(pltxack), .b(net11), .c(net30) );
    oa21_1 \U149/U1  ( .x(\U149/n2 ), .a(\U149/n2 ), .b(\U149/nr ), .c(
        \U149/nd ) );
    inv_2 \U149/U3  ( .x(txdone), .a(\U149/n2 ) );
    inv_1 \U133/U618/U3  ( .x(net23), .a(net15) );
    inv_1 \U133/U617/U3  ( .x(net25), .a(routetxreq) );
    ao23_1 \U133/U616/U21/U1/U1  ( .x(routetxreq), .a(pltxreq), .b(routetxreq), 
        .c(pltxreq), .d(\locked[0] ), .e(net23) );
    ao23_1 \U133/U615/U21/U1/U1  ( .x(net15), .a(pltxreq), .b(net15), .c(
        pltxreq), .d(\locked[1] ), .e(net25) );
    and2_1 \U160/U2/U8  ( .x(lwrite), .a(candefer), .b(\U160/acb ) );
    nor2_1 \U160/U3/U5  ( .x(net30), .a(\U160/acb ), .b(net26) );
    oai21_1 \U160/U1/U30/U1/U1  ( .x(\U160/acb ), .a(\U160/U1/Z ), .b(net26), 
        .c(candefer) );
    inv_1 \U160/U1/U30/U1/U2  ( .x(\U160/U1/Z ), .a(\U160/acb ) );
    nand3_2 \U136/U48/U16  ( .x(\locked[0] ), .a(\locked[1] ), .b(
        \U136/nclear_latch ), .c(\U136/nwl ) );
    nor2_0 \U136/U36/U5  ( .x(\U136/nulsense ), .a(\locked[1] ), .b(\U136/nwl 
        ) );
    nor2_0 \U136/U37/U5  ( .x(\U136/nlsense ), .a(\U136/nwh ), .b(\locked[0] )
         );
    and2_1 \U136/U76/U8  ( .x(\U136/nclear_latch ), .a(nReset), .b(nlclear) );
    nor2_1 \U136/U77/U5  ( .x(lockcleared), .a(nlclear), .b(\locked[1] ) );
    nand2_1 \U136/U14/U5  ( .x(\U136/nwl ), .a(lwrite), .b(n2) );
    nand2_1 \U136/U15/U5  ( .x(\U136/nwh ), .a(n1), .b(lwrite) );
    nand2_2 \U136/U47/U5  ( .x(\locked[1] ), .a(\U136/nwh ), .b(\locked[0] )
         );
    or2_4 \U136/U35/U12  ( .x(net26), .a(\U136/nlsense ), .b(\U136/nulsense )
         );
    buf_1 U1 ( .x(n1), .a(lock[1]) );
    buf_1 U2 ( .x(n2), .a(lock[0]) );
endmodule


module chain_irdemuxNew_1 ( err, ncback, rd, rnw, status, cbh, cbl, nReset, 
    nack, statusack );
output [1:0] err;
output [63:0] rd;
output [1:0] rnw;
output [1:0] status;
input  [7:0] cbh;
input  [7:0] cbl;
input  nReset, nack, statusack;
output ncback;
    wire n17, n18, \ncd[7] , \ncd[6] , \ncd[5] , \ncd[4] , \ncd[3] , \ncd[2] , 
        \ncd[1] , \ncd[0] , \col_h[2] , \col_h[1] , \col_h[0] , \col_l[2] , 
        \col_l[1] , \col_l[0] , \opc_l[2] , \opc_l[1] , \opc_l[0] , \opc_h[1] , 
        \opc_h[0] , pullcd, net86, net171, net168, net103, net170, bpullcd, 
        reset, net94, read_lhw, net166, net169, read, net139, net172, 
        start_receiving, net193, net167, net149, net173, pkt_normal, notify, 
        net150, write, net176, net162, pkt_done, net0187, net0208, 
        \U1697/U21/nr , \U1697/U21/nd , \U1697/U21/n2 , \U307/U21/nr , 
        \U307/U21/nd , \U307/U21/n2 , \U1664/U28/Z , \U1664/U32/Z , 
        \U1664/U29/Z , \U1664/U33/Z , \U1664/U30/Z , \U1664/U31/Z , 
        \U1664/U37/Z , \U1664/y[0] , \U1664/y[1] , \U1664/x[1] , \U1664/x[3] , 
        \U1664/x[2] , \U1664/x[0] , \U1698/nr , \U1698/nd , \U1698/n2 , 
        \I6/oh[7] , \I6/oh[6] , \I6/oh[4] , \I6/oh[3] , \I6/oh[2] , \I6/ol[7] , 
        \I6/ol[6] , \I6/ol[4] , \I6/ol[3] , \I6/drivel , \I6/driveh , 
        \I6/localcd , \I6/ncd[7] , \I6/ncd[6] , \I6/ncd[5] , \I6/ncd[4] , 
        \I6/ncd[3] , \I6/ncd[2] , \I6/ncd[1] , \I6/ncd[0] , \I6/ba , 
        \I6/latch , \I6/acb , \I6/ctrlack_internal , \I6/nlocalcd , 
        \I6/U4/U28/U1/clr , \I6/U4/U28/U1/set , \I6/U1/Z , \I6/U1664/y[0] , 
        \I6/U1664/y[1] , \I6/U1664/x[1] , \I6/U1664/x[3] , \I6/U1664/x[2] , 
        \I6/U1664/x[0] , \I6/U1664/U28/Z , \I6/U1664/U32/Z , \I6/U1664/U29/Z , 
        \I6/U1664/U33/Z , \I6/U1664/U30/Z , \I6/U1664/U31/Z , \I6/U1664/U37/Z , 
        \I6/U1669/nr , \I6/U1669/nd , \I6/U1669/n2 , \U1667/drivel , 
        \U1667/driveh , \U1667/localcd , \U1667/ncd[7] , \U1667/ncd[6] , 
        \U1667/ncd[5] , \U1667/ncd[4] , \U1667/ncd[3] , \U1667/ncd[2] , 
        \U1667/ncd[1] , \U1667/ncd[0] , \U1667/ba , \U1667/latch , \U1667/acb , 
        \U1667/ctrlack_internal , \U1667/nlocalcd , \U1667/U4/U28/U1/clr , 
        \U1667/U4/U28/U1/set , \U1667/U1/Z , \U1667/U1664/y[0] , 
        \U1667/U1664/y[1] , \U1667/U1664/x[1] , \U1667/U1664/x[3] , 
        \U1667/U1664/x[2] , \U1667/U1664/x[0] , \U1667/U1664/U28/Z , 
        \U1667/U1664/U32/Z , \U1667/U1664/U29/Z , \U1667/U1664/U33/Z , 
        \U1667/U1664/U30/Z , \U1667/U1664/U31/Z , \U1667/U1664/U37/Z , 
        \U1667/U1669/nr , \U1667/U1669/nd , \U1667/U1669/n2 , \U1650/oh[4] , 
        \U1650/oh[3] , \U1650/oh[2] , \U1650/oh[1] , \U1650/oh[0] , 
        \U1650/ol[4] , \U1650/ol[3] , \U1650/ol[2] , \U1650/ol[1] , 
        \U1650/ol[0] , \U1650/drivel , \U1650/driveh , \U1650/localcd , 
        \U1650/ncd[7] , \U1650/ncd[6] , \U1650/ncd[5] , \U1650/ncd[4] , 
        \U1650/ncd[3] , \U1650/ncd[2] , \U1650/ncd[1] , \U1650/ncd[0] , 
        \U1650/ba , \U1650/latch , \U1650/acb , \U1650/ctrlack_internal , 
        \U1650/nlocalcd , \U1650/U4/U28/U1/clr , \U1650/U4/U28/U1/set , 
        \U1650/U1/Z , \U1650/U1664/y[0] , \U1650/U1664/y[1] , 
        \U1650/U1664/x[1] , \U1650/U1664/x[3] , \U1650/U1664/x[2] , 
        \U1650/U1664/x[0] , \U1650/U1664/U28/Z , \U1650/U1664/U32/Z , 
        \U1650/U1664/U29/Z , \U1650/U1664/U33/Z , \U1650/U1664/U30/Z , 
        \U1650/U1664/U31/Z , \U1650/U1664/U37/Z , \U1650/U1669/nr , 
        \U1650/U1669/nd , \U1650/U1669/n2 , \U1666/drivel , \U1666/driveh , 
        \U1666/localcd , \U1666/ncd[7] , \U1666/ncd[6] , \U1666/ncd[5] , 
        \U1666/ncd[4] , \U1666/ncd[3] , \U1666/ncd[2] , \U1666/ncd[1] , 
        \U1666/ncd[0] , \U1666/ba , \U1666/latch , \U1666/acb , 
        \U1666/ctrlack_internal , \U1666/nlocalcd , \U1666/U4/U28/U1/clr , 
        \U1666/U4/U28/U1/set , \U1666/U1/Z , \U1666/U1664/y[0] , 
        \U1666/U1664/y[1] , \U1666/U1664/x[1] , \U1666/U1664/x[3] , 
        \U1666/U1664/x[2] , \U1666/U1664/x[0] , \U1666/U1664/U28/Z , 
        \U1666/U1664/U32/Z , \U1666/U1664/U29/Z , \U1666/U1664/U33/Z , 
        \U1666/U1664/U30/Z , \U1666/U1664/U31/Z , \U1666/U1664/U37/Z , 
        \U1666/U1669/nr , \U1666/U1669/nd , \U1666/U1669/n2 , \I1/drivel , 
        \I1/driveh , \I1/localcd , \I1/ncd[7] , \I1/ncd[6] , \I1/ncd[5] , 
        \I1/ncd[4] , \I1/ncd[3] , \I1/ncd[2] , \I1/ncd[1] , \I1/ncd[0] , 
        \I1/ba , \I1/latch , \I1/acb , \I1/ctrlack_internal , \I1/nlocalcd , 
        \I1/U4/U28/U1/clr , \I1/U4/U28/U1/set , \I1/U1/Z , \I1/U1664/y[0] , 
        \I1/U1664/y[1] , \I1/U1664/x[1] , \I1/U1664/x[3] , \I1/U1664/x[2] , 
        \I1/U1664/x[0] , \I1/U1664/U28/Z , \I1/U1664/U32/Z , \I1/U1664/U29/Z , 
        \I1/U1664/U33/Z , \I1/U1664/U30/Z , \I1/U1664/U31/Z , \I1/U1664/U37/Z , 
        \I1/U1669/nr , \I1/U1669/nd , \I1/U1669/n2 , \I2/drivel , \I2/driveh , 
        \I2/localcd , \I2/ncd[7] , \I2/ncd[6] , \I2/ncd[5] , \I2/ncd[4] , 
        \I2/ncd[3] , \I2/ncd[2] , \I2/ncd[1] , \I2/ncd[0] , \I2/ba , 
        \I2/latch , \I2/acb , \I2/ctrlack_internal , \I2/nlocalcd , 
        \I2/U4/U28/U1/clr , \I2/U4/U28/U1/set , \I2/U1/Z , \I2/U1664/y[0] , 
        \I2/U1664/y[1] , \I2/U1664/x[1] , \I2/U1664/x[3] , \I2/U1664/x[2] , 
        \I2/U1664/x[0] , \I2/U1664/U28/Z , \I2/U1664/U32/Z , \I2/U1664/U29/Z , 
        \I2/U1664/U33/Z , \I2/U1664/U30/Z , \I2/U1664/U31/Z , \I2/U1664/U37/Z , 
        \I2/U1669/nr , \I2/U1669/nd , \I2/U1669/n2 , n1, n2, n3, n4, n5, n6, 
        n7, n8, n9, n10, n11, n12, n13, n14;
    buf_1 U262 ( .x(bpullcd), .a(pullcd) );
    or2_4 \U1674/U12  ( .x(net162), .a(nack), .b(reset) );
    and2_4 \U1785/U8  ( .x(pkt_normal), .a(\opc_l[2] ), .b(\opc_l[1] ) );
    and2_4 \U1777/U8  ( .x(net150), .a(\opc_l[2] ), .b(\opc_h[1] ) );
    or3_1 \U1813/U12  ( .x(pkt_done), .a(write), .b(reset), .c(net193) );
    nor2_1 \U1651_0_/U5  ( .x(\ncd[0] ), .a(cbh[0]), .b(cbl[0]) );
    nor2_1 \U1651_1_/U5  ( .x(\ncd[1] ), .a(cbh[1]), .b(cbl[1]) );
    nor2_1 \U1651_2_/U5  ( .x(\ncd[2] ), .a(cbh[2]), .b(cbl[2]) );
    nor2_1 \U1651_3_/U5  ( .x(\ncd[3] ), .a(cbh[3]), .b(cbl[3]) );
    nor2_1 \U1651_4_/U5  ( .x(\ncd[4] ), .a(cbh[4]), .b(cbl[4]) );
    nor2_1 \U1651_5_/U5  ( .x(\ncd[5] ), .a(cbh[5]), .b(cbl[5]) );
    nor2_1 \U1651_6_/U5  ( .x(\ncd[6] ), .a(cbh[6]), .b(cbl[6]) );
    nor2_1 \U1651_7_/U5  ( .x(\ncd[7] ), .a(cbh[7]), .b(cbl[7]) );
    nor2_1 \U1812/U5  ( .x(start_receiving), .a(notify), .b(net176) );
    nor2_1 \I7/U5  ( .x(net86), .a(net172), .b(net173) );
    nor2_1 \I4/U5  ( .x(net171), .a(net169), .b(net170) );
    nor2_1 \I3/U5  ( .x(net168), .a(net166), .b(net167) );
    inv_2 \U1675/U3  ( .x(reset), .a(nReset) );
    nand3_2 \U193/U16  ( .x(ncback), .a(net86), .b(net171), .c(net168) );
    ao222_1 \U1811/U18/U1/U1  ( .x(net176), .a(net162), .b(pkt_done), .c(
        net162), .d(net176), .e(pkt_done), .f(net176) );
    aoi222_1 \U1664/U28/U30/U1  ( .x(\U1664/x[3] ), .a(\ncd[7] ), .b(\ncd[6] ), 
        .c(\ncd[7] ), .d(\U1664/U28/Z ), .e(\ncd[6] ), .f(\U1664/U28/Z ) );
    inv_1 \U1664/U28/U30/Uinv  ( .x(\U1664/U28/Z ), .a(\U1664/x[3] ) );
    aoi222_1 \U1664/U32/U30/U1  ( .x(\U1664/x[0] ), .a(\ncd[1] ), .b(\ncd[0] ), 
        .c(\ncd[1] ), .d(\U1664/U32/Z ), .e(\ncd[0] ), .f(\U1664/U32/Z ) );
    inv_1 \U1664/U32/U30/Uinv  ( .x(\U1664/U32/Z ), .a(\U1664/x[0] ) );
    aoi222_1 \U1664/U29/U30/U1  ( .x(\U1664/x[2] ), .a(\ncd[5] ), .b(\ncd[4] ), 
        .c(\ncd[5] ), .d(\U1664/U29/Z ), .e(\ncd[4] ), .f(\U1664/U29/Z ) );
    inv_1 \U1664/U29/U30/Uinv  ( .x(\U1664/U29/Z ), .a(\U1664/x[2] ) );
    aoi222_1 \U1664/U33/U30/U1  ( .x(\U1664/y[0] ), .a(\U1664/x[1] ), .b(
        \U1664/x[0] ), .c(\U1664/x[1] ), .d(\U1664/U33/Z ), .e(\U1664/x[0] ), 
        .f(\U1664/U33/Z ) );
    inv_1 \U1664/U33/U30/Uinv  ( .x(\U1664/U33/Z ), .a(\U1664/y[0] ) );
    aoi222_1 \U1664/U30/U30/U1  ( .x(\U1664/y[1] ), .a(\U1664/x[3] ), .b(
        \U1664/x[2] ), .c(\U1664/x[3] ), .d(\U1664/U30/Z ), .e(\U1664/x[2] ), 
        .f(\U1664/U30/Z ) );
    inv_1 \U1664/U30/U30/Uinv  ( .x(\U1664/U30/Z ), .a(\U1664/y[1] ) );
    aoi222_1 \U1664/U31/U30/U1  ( .x(\U1664/x[1] ), .a(\ncd[3] ), .b(\ncd[2] ), 
        .c(\ncd[3] ), .d(\U1664/U31/Z ), .e(\ncd[2] ), .f(\U1664/U31/Z ) );
    inv_1 \U1664/U31/U30/Uinv  ( .x(\U1664/U31/Z ), .a(\U1664/x[1] ) );
    aoi222_1 \U1664/U37/U30/U1  ( .x(pullcd), .a(\U1664/y[0] ), .b(
        \U1664/y[1] ), .c(\U1664/y[0] ), .d(\U1664/U37/Z ), .e(\U1664/y[1] ), 
        .f(\U1664/U37/Z ) );
    inv_1 \U1664/U37/U30/Uinv  ( .x(\U1664/U37/Z ), .a(pullcd) );
    nor3_1 \U1697/U21/Unr  ( .x(\U1697/U21/nr ), .a(rnw[0]), .b(pkt_normal), 
        .c(net149) );
    nand3_1 \U1697/U21/Und  ( .x(\U1697/U21/nd ), .a(rnw[0]), .b(pkt_normal), 
        .c(net149) );
    oa21_1 \U1697/U21/U1  ( .x(\U1697/U21/n2 ), .a(\U1697/U21/n2 ), .b(
        \U1697/U21/nr ), .c(\U1697/U21/nd ) );
    inv_1 \U1697/U21/U3  ( .x(write), .a(\U1697/U21/n2 ) );
    nor3_1 \U307/U21/Unr  ( .x(\U307/U21/nr ), .a(net149), .b(net150), .c(
        statusack) );
    nand3_1 \U307/U21/Und  ( .x(\U307/U21/nd ), .a(net149), .b(net150), .c(
        statusack) );
    oa21_1 \U307/U21/U1  ( .x(\U307/U21/n2 ), .a(\U307/U21/n2 ), .b(
        \U307/U21/nr ), .c(\U307/U21/nd ) );
    inv_1 \U307/U21/U3  ( .x(notify), .a(\U307/U21/n2 ) );
    nor3_1 \U1698/Unr  ( .x(\U1698/nr ), .a(rnw[1]), .b(pkt_normal), .c(net149
        ) );
    nand3_1 \U1698/Und  ( .x(\U1698/nd ), .a(rnw[1]), .b(pkt_normal), .c(
        net149) );
    oa21_1 \U1698/U1  ( .x(\U1698/n2 ), .a(\U1698/n2 ), .b(\U1698/nr ), .c(
        \U1698/nd ) );
    inv_2 \U1698/U3  ( .x(read), .a(\U1698/n2 ) );
    and2_1 \U1756/U1754/U8  ( .x(n17), .a(\opc_h[0] ), .b(pkt_normal) );
    and2_1 \U1756/U1755/U8  ( .x(n18), .a(\opc_l[0] ), .b(pkt_normal) );
    and2_1 \U1800/U1754/U8  ( .x(rnw[1]), .a(net0187), .b(pkt_normal) );
    and2_1 \U1800/U1755/U8  ( .x(rnw[0]), .a(net0208), .b(pkt_normal) );
    and2_1 \U1758/U1754/U8  ( .x(status[1]), .a(\opc_h[0] ), .b(net150) );
    and2_1 \U1758/U1755/U8  ( .x(status[0]), .a(\opc_l[0] ), .b(net150) );
    buf_2 \I6/U1653  ( .x(\I6/latch ), .a(net173) );
    nor2_1 \I6/U264/U5  ( .x(\I6/nlocalcd ), .a(reset), .b(\I6/localcd ) );
    nor2_1 \I6/U1659_0_/U5  ( .x(\I6/ncd[0] ), .a(\opc_l[0] ), .b(\opc_h[0] )
         );
    nor2_1 \I6/U1659_1_/U5  ( .x(\I6/ncd[1] ), .a(\opc_l[1] ), .b(\opc_h[1] )
         );
    nor2_1 \I6/U1659_2_/U5  ( .x(\I6/ncd[2] ), .a(\opc_l[2] ), .b(\I6/oh[2] )
         );
    nor2_1 \I6/U1659_3_/U5  ( .x(\I6/ncd[3] ), .a(\I6/ol[3] ), .b(\I6/oh[3] )
         );
    nor2_1 \I6/U1659_4_/U5  ( .x(\I6/ncd[4] ), .a(\I6/ol[4] ), .b(\I6/oh[4] )
         );
    nor2_1 \I6/U1659_5_/U5  ( .x(\I6/ncd[5] ), .a(net0208), .b(net0187) );
    nor2_1 \I6/U1659_6_/U5  ( .x(\I6/ncd[6] ), .a(\I6/ol[6] ), .b(\I6/oh[6] )
         );
    nor2_1 \I6/U1659_7_/U5  ( .x(\I6/ncd[7] ), .a(\I6/ol[7] ), .b(\I6/oh[7] )
         );
    nor2_1 \I6/U3/U5  ( .x(\I6/ctrlack_internal ), .a(\I6/acb ), .b(\I6/ba )
         );
    buf_2 \I6/U1665/U7  ( .x(\I6/driveh ), .a(net139) );
    buf_2 \I6/U1666/U7  ( .x(\I6/drivel ), .a(net139) );
    ao23_1 \I6/U1658_0_/U21/U1/U1  ( .x(\opc_l[0] ), .a(\I6/driveh ), .b(
        \opc_l[0] ), .c(\I6/driveh ), .d(cbl[0]), .e(n12) );
    ao23_1 \I6/U1658_1_/U21/U1/U1  ( .x(\opc_l[1] ), .a(\I6/driveh ), .b(
        \opc_l[1] ), .c(\I6/drivel ), .d(cbl[1]), .e(n12) );
    ao23_1 \I6/U1658_2_/U21/U1/U1  ( .x(\opc_l[2] ), .a(\I6/drivel ), .b(
        \opc_l[2] ), .c(n13), .d(cbl[2]), .e(n12) );
    ao23_1 \I6/U1658_3_/U21/U1/U1  ( .x(\I6/ol[3] ), .a(\I6/drivel ), .b(
        \I6/ol[3] ), .c(\I6/drivel ), .d(cbl[3]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_4_/U21/U1/U1  ( .x(\I6/ol[4] ), .a(n13), .b(\I6/ol[4] ), 
        .c(n13), .d(cbl[4]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_5_/U21/U1/U1  ( .x(net0208), .a(\I6/driveh ), .b(net0208), 
        .c(\I6/driveh ), .d(cbl[5]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_6_/U21/U1/U1  ( .x(\I6/ol[6] ), .a(n13), .b(\I6/ol[6] ), 
        .c(n13), .d(cbl[6]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_7_/U21/U1/U1  ( .x(\I6/ol[7] ), .a(n13), .b(\I6/ol[7] ), 
        .c(\I6/driveh ), .d(cbl[7]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_0_/U21/U1/U1  ( .x(\opc_h[0] ), .a(n13), .b(\opc_h[0] ), 
        .c(\I6/drivel ), .d(cbh[0]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_1_/U21/U1/U1  ( .x(\opc_h[1] ), .a(\I6/driveh ), .b(
        \opc_h[1] ), .c(n13), .d(cbh[1]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_2_/U21/U1/U1  ( .x(\I6/oh[2] ), .a(\I6/driveh ), .b(
        \I6/oh[2] ), .c(n13), .d(cbh[2]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_3_/U21/U1/U1  ( .x(\I6/oh[3] ), .a(\I6/drivel ), .b(
        \I6/oh[3] ), .c(\I6/drivel ), .d(cbh[3]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_4_/U21/U1/U1  ( .x(\I6/oh[4] ), .a(n13), .b(\I6/oh[4] ), 
        .c(\I6/driveh ), .d(cbh[4]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_5_/U21/U1/U1  ( .x(net0187), .a(\I6/driveh ), .b(net0187), 
        .c(\I6/driveh ), .d(cbh[5]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_6_/U21/U1/U1  ( .x(\I6/oh[6] ), .a(\I6/drivel ), .b(
        \I6/oh[6] ), .c(\I6/drivel ), .d(cbh[6]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_7_/U21/U1/U1  ( .x(\I6/oh[7] ), .a(\I6/drivel ), .b(
        \I6/oh[7] ), .c(n13), .d(cbh[7]), .e(\I6/latch ) );
    aoai211_1 \I6/U4/U28/U1/U1  ( .x(\I6/U4/U28/U1/clr ), .a(net139), .b(
        \I6/acb ), .c(\I6/nlocalcd ), .d(net173) );
    nand3_1 \I6/U4/U28/U1/U2  ( .x(\I6/U4/U28/U1/set ), .a(\I6/nlocalcd ), .b(
        net139), .c(\I6/acb ) );
    nand2_2 \I6/U4/U28/U1/U3  ( .x(net173), .a(\I6/U4/U28/U1/clr ), .b(
        \I6/U4/U28/U1/set ) );
    oai21_1 \I6/U1/U30/U1/U1  ( .x(\I6/acb ), .a(\I6/U1/Z ), .b(\I6/ba ), .c(
        net139) );
    inv_1 \I6/U1/U30/U1/U2  ( .x(\I6/U1/Z ), .a(\I6/acb ) );
    ao222_1 \I6/U5/U18/U1/U1  ( .x(\I6/ba ), .a(\I6/latch ), .b(n14), .c(
        \I6/latch ), .d(\I6/ba ), .e(n14), .f(\I6/ba ) );
    aoi222_1 \I6/U1664/U28/U30/U1  ( .x(\I6/U1664/x[3] ), .a(\I6/ncd[7] ), .b(
        \I6/ncd[6] ), .c(\I6/ncd[7] ), .d(\I6/U1664/U28/Z ), .e(\I6/ncd[6] ), 
        .f(\I6/U1664/U28/Z ) );
    inv_1 \I6/U1664/U28/U30/Uinv  ( .x(\I6/U1664/U28/Z ), .a(\I6/U1664/x[3] )
         );
    aoi222_1 \I6/U1664/U32/U30/U1  ( .x(\I6/U1664/x[0] ), .a(\I6/ncd[1] ), .b(
        \I6/ncd[0] ), .c(\I6/ncd[1] ), .d(\I6/U1664/U32/Z ), .e(\I6/ncd[0] ), 
        .f(\I6/U1664/U32/Z ) );
    inv_1 \I6/U1664/U32/U30/Uinv  ( .x(\I6/U1664/U32/Z ), .a(\I6/U1664/x[0] )
         );
    aoi222_1 \I6/U1664/U29/U30/U1  ( .x(\I6/U1664/x[2] ), .a(\I6/ncd[5] ), .b(
        \I6/ncd[4] ), .c(\I6/ncd[5] ), .d(\I6/U1664/U29/Z ), .e(\I6/ncd[4] ), 
        .f(\I6/U1664/U29/Z ) );
    inv_1 \I6/U1664/U29/U30/Uinv  ( .x(\I6/U1664/U29/Z ), .a(\I6/U1664/x[2] )
         );
    aoi222_1 \I6/U1664/U33/U30/U1  ( .x(\I6/U1664/y[0] ), .a(\I6/U1664/x[1] ), 
        .b(\I6/U1664/x[0] ), .c(\I6/U1664/x[1] ), .d(\I6/U1664/U33/Z ), .e(
        \I6/U1664/x[0] ), .f(\I6/U1664/U33/Z ) );
    inv_1 \I6/U1664/U33/U30/Uinv  ( .x(\I6/U1664/U33/Z ), .a(\I6/U1664/y[0] )
         );
    aoi222_1 \I6/U1664/U30/U30/U1  ( .x(\I6/U1664/y[1] ), .a(\I6/U1664/x[3] ), 
        .b(\I6/U1664/x[2] ), .c(\I6/U1664/x[3] ), .d(\I6/U1664/U30/Z ), .e(
        \I6/U1664/x[2] ), .f(\I6/U1664/U30/Z ) );
    inv_1 \I6/U1664/U30/U30/Uinv  ( .x(\I6/U1664/U30/Z ), .a(\I6/U1664/y[1] )
         );
    aoi222_1 \I6/U1664/U31/U30/U1  ( .x(\I6/U1664/x[1] ), .a(\I6/ncd[3] ), .b(
        \I6/ncd[2] ), .c(\I6/ncd[3] ), .d(\I6/U1664/U31/Z ), .e(\I6/ncd[2] ), 
        .f(\I6/U1664/U31/Z ) );
    inv_1 \I6/U1664/U31/U30/Uinv  ( .x(\I6/U1664/U31/Z ), .a(\I6/U1664/x[1] )
         );
    aoi222_1 \I6/U1664/U37/U30/U1  ( .x(\I6/localcd ), .a(\I6/U1664/y[0] ), 
        .b(\I6/U1664/y[1] ), .c(\I6/U1664/y[0] ), .d(\I6/U1664/U37/Z ), .e(
        \I6/U1664/y[1] ), .f(\I6/U1664/U37/Z ) );
    inv_1 \I6/U1664/U37/U30/Uinv  ( .x(\I6/U1664/U37/Z ), .a(\I6/localcd ) );
    nor3_1 \I6/U1669/Unr  ( .x(\I6/U1669/nr ), .a(\I6/ctrlack_internal ), .b(
        n13), .c(\I6/drivel ) );
    nand3_1 \I6/U1669/Und  ( .x(\I6/U1669/nd ), .a(\I6/ctrlack_internal ), .b(
        \I6/driveh ), .c(\I6/drivel ) );
    oa21_1 \I6/U1669/U1  ( .x(\I6/U1669/n2 ), .a(\I6/U1669/n2 ), .b(
        \I6/U1669/nr ), .c(\I6/U1669/nd ) );
    inv_2 \I6/U1669/U3  ( .x(net149), .a(\I6/U1669/n2 ) );
    buf_2 \U1667/U1653  ( .x(\U1667/latch ), .a(net167) );
    nor2_1 \U1667/U264/U5  ( .x(\U1667/nlocalcd ), .a(reset), .b(
        \U1667/localcd ) );
    nor2_1 \U1667/U1659_0_/U5  ( .x(\U1667/ncd[0] ), .a(rd[0]), .b(rd[32]) );
    nor2_1 \U1667/U1659_1_/U5  ( .x(\U1667/ncd[1] ), .a(rd[1]), .b(rd[33]) );
    nor2_1 \U1667/U1659_2_/U5  ( .x(\U1667/ncd[2] ), .a(rd[2]), .b(rd[34]) );
    nor2_1 \U1667/U1659_3_/U5  ( .x(\U1667/ncd[3] ), .a(rd[3]), .b(rd[35]) );
    nor2_1 \U1667/U1659_4_/U5  ( .x(\U1667/ncd[4] ), .a(rd[4]), .b(rd[36]) );
    nor2_1 \U1667/U1659_5_/U5  ( .x(\U1667/ncd[5] ), .a(rd[5]), .b(rd[37]) );
    nor2_1 \U1667/U1659_6_/U5  ( .x(\U1667/ncd[6] ), .a(rd[6]), .b(rd[38]) );
    nor2_1 \U1667/U1659_7_/U5  ( .x(\U1667/ncd[7] ), .a(rd[7]), .b(rd[39]) );
    nor2_1 \U1667/U3/U5  ( .x(\U1667/ctrlack_internal ), .a(\U1667/acb ), .b(
        \U1667/ba ) );
    buf_2 \U1667/U1665/U7  ( .x(\U1667/driveh ), .a(read_lhw) );
    buf_2 \U1667/U1666/U7  ( .x(\U1667/drivel ), .a(read_lhw) );
    ao23_1 \U1667/U1658_0_/U21/U1/U1  ( .x(rd[0]), .a(n11), .b(rd[0]), .c(
        \U1667/drivel ), .d(cbl[0]), .e(n10) );
    ao23_1 \U1667/U1658_1_/U21/U1/U1  ( .x(rd[1]), .a(n11), .b(rd[1]), .c(
        \U1667/driveh ), .d(cbl[1]), .e(n10) );
    ao23_1 \U1667/U1658_2_/U21/U1/U1  ( .x(rd[2]), .a(\U1667/driveh ), .b(rd
        [2]), .c(n11), .d(cbl[2]), .e(n10) );
    ao23_1 \U1667/U1658_3_/U21/U1/U1  ( .x(rd[3]), .a(n11), .b(rd[3]), .c(
        \U1667/driveh ), .d(cbl[3]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_4_/U21/U1/U1  ( .x(rd[4]), .a(\U1667/drivel ), .b(rd
        [4]), .c(n11), .d(cbl[4]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_5_/U21/U1/U1  ( .x(rd[5]), .a(\U1667/drivel ), .b(rd
        [5]), .c(n11), .d(cbl[5]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_6_/U21/U1/U1  ( .x(rd[6]), .a(\U1667/driveh ), .b(rd
        [6]), .c(\U1667/drivel ), .d(cbl[6]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_7_/U21/U1/U1  ( .x(rd[7]), .a(\U1667/driveh ), .b(rd
        [7]), .c(\U1667/driveh ), .d(cbl[7]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_0_/U21/U1/U1  ( .x(rd[32]), .a(\U1667/drivel ), .b(rd
        [32]), .c(n11), .d(cbh[0]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_1_/U21/U1/U1  ( .x(rd[33]), .a(\U1667/driveh ), .b(rd
        [33]), .c(\U1667/drivel ), .d(cbh[1]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_2_/U21/U1/U1  ( .x(rd[34]), .a(\U1667/drivel ), .b(rd
        [34]), .c(\U1667/drivel ), .d(cbh[2]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_3_/U21/U1/U1  ( .x(rd[35]), .a(\U1667/driveh ), .b(rd
        [35]), .c(\U1667/driveh ), .d(cbh[3]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_4_/U21/U1/U1  ( .x(rd[36]), .a(\U1667/drivel ), .b(rd
        [36]), .c(\U1667/driveh ), .d(cbh[4]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_5_/U21/U1/U1  ( .x(rd[37]), .a(\U1667/driveh ), .b(rd
        [37]), .c(n11), .d(cbh[5]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_6_/U21/U1/U1  ( .x(rd[38]), .a(n11), .b(rd[38]), .c(
        \U1667/drivel ), .d(cbh[6]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_7_/U21/U1/U1  ( .x(rd[39]), .a(n11), .b(rd[39]), .c(
        n11), .d(cbh[7]), .e(\U1667/latch ) );
    aoai211_1 \U1667/U4/U28/U1/U1  ( .x(\U1667/U4/U28/U1/clr ), .a(read_lhw), 
        .b(\U1667/acb ), .c(\U1667/nlocalcd ), .d(net167) );
    nand3_1 \U1667/U4/U28/U1/U2  ( .x(\U1667/U4/U28/U1/set ), .a(
        \U1667/nlocalcd ), .b(read_lhw), .c(\U1667/acb ) );
    nand2_2 \U1667/U4/U28/U1/U3  ( .x(net167), .a(\U1667/U4/U28/U1/clr ), .b(
        \U1667/U4/U28/U1/set ) );
    oai21_1 \U1667/U1/U30/U1/U1  ( .x(\U1667/acb ), .a(\U1667/U1/Z ), .b(
        \U1667/ba ), .c(read_lhw) );
    inv_1 \U1667/U1/U30/U1/U2  ( .x(\U1667/U1/Z ), .a(\U1667/acb ) );
    ao222_1 \U1667/U5/U18/U1/U1  ( .x(\U1667/ba ), .a(\U1667/latch ), .b(n14), 
        .c(\U1667/latch ), .d(\U1667/ba ), .e(n14), .f(\U1667/ba ) );
    aoi222_1 \U1667/U1664/U28/U30/U1  ( .x(\U1667/U1664/x[3] ), .a(
        \U1667/ncd[7] ), .b(\U1667/ncd[6] ), .c(\U1667/ncd[7] ), .d(
        \U1667/U1664/U28/Z ), .e(\U1667/ncd[6] ), .f(\U1667/U1664/U28/Z ) );
    inv_1 \U1667/U1664/U28/U30/Uinv  ( .x(\U1667/U1664/U28/Z ), .a(
        \U1667/U1664/x[3] ) );
    aoi222_1 \U1667/U1664/U32/U30/U1  ( .x(\U1667/U1664/x[0] ), .a(
        \U1667/ncd[1] ), .b(\U1667/ncd[0] ), .c(\U1667/ncd[1] ), .d(
        \U1667/U1664/U32/Z ), .e(\U1667/ncd[0] ), .f(\U1667/U1664/U32/Z ) );
    inv_1 \U1667/U1664/U32/U30/Uinv  ( .x(\U1667/U1664/U32/Z ), .a(
        \U1667/U1664/x[0] ) );
    aoi222_1 \U1667/U1664/U29/U30/U1  ( .x(\U1667/U1664/x[2] ), .a(
        \U1667/ncd[5] ), .b(\U1667/ncd[4] ), .c(\U1667/ncd[5] ), .d(
        \U1667/U1664/U29/Z ), .e(\U1667/ncd[4] ), .f(\U1667/U1664/U29/Z ) );
    inv_1 \U1667/U1664/U29/U30/Uinv  ( .x(\U1667/U1664/U29/Z ), .a(
        \U1667/U1664/x[2] ) );
    aoi222_1 \U1667/U1664/U33/U30/U1  ( .x(\U1667/U1664/y[0] ), .a(
        \U1667/U1664/x[1] ), .b(\U1667/U1664/x[0] ), .c(\U1667/U1664/x[1] ), 
        .d(\U1667/U1664/U33/Z ), .e(\U1667/U1664/x[0] ), .f(
        \U1667/U1664/U33/Z ) );
    inv_1 \U1667/U1664/U33/U30/Uinv  ( .x(\U1667/U1664/U33/Z ), .a(
        \U1667/U1664/y[0] ) );
    aoi222_1 \U1667/U1664/U30/U30/U1  ( .x(\U1667/U1664/y[1] ), .a(
        \U1667/U1664/x[3] ), .b(\U1667/U1664/x[2] ), .c(\U1667/U1664/x[3] ), 
        .d(\U1667/U1664/U30/Z ), .e(\U1667/U1664/x[2] ), .f(
        \U1667/U1664/U30/Z ) );
    inv_1 \U1667/U1664/U30/U30/Uinv  ( .x(\U1667/U1664/U30/Z ), .a(
        \U1667/U1664/y[1] ) );
    aoi222_1 \U1667/U1664/U31/U30/U1  ( .x(\U1667/U1664/x[1] ), .a(
        \U1667/ncd[3] ), .b(\U1667/ncd[2] ), .c(\U1667/ncd[3] ), .d(
        \U1667/U1664/U31/Z ), .e(\U1667/ncd[2] ), .f(\U1667/U1664/U31/Z ) );
    inv_1 \U1667/U1664/U31/U30/Uinv  ( .x(\U1667/U1664/U31/Z ), .a(
        \U1667/U1664/x[1] ) );
    aoi222_1 \U1667/U1664/U37/U30/U1  ( .x(\U1667/localcd ), .a(
        \U1667/U1664/y[0] ), .b(\U1667/U1664/y[1] ), .c(\U1667/U1664/y[0] ), 
        .d(\U1667/U1664/U37/Z ), .e(\U1667/U1664/y[1] ), .f(
        \U1667/U1664/U37/Z ) );
    inv_1 \U1667/U1664/U37/U30/Uinv  ( .x(\U1667/U1664/U37/Z ), .a(
        \U1667/localcd ) );
    nor3_1 \U1667/U1669/Unr  ( .x(\U1667/U1669/nr ), .a(
        \U1667/ctrlack_internal ), .b(n11), .c(\U1667/drivel ) );
    nand3_1 \U1667/U1669/Und  ( .x(\U1667/U1669/nd ), .a(
        \U1667/ctrlack_internal ), .b(\U1667/driveh ), .c(\U1667/drivel ) );
    oa21_1 \U1667/U1669/U1  ( .x(\U1667/U1669/n2 ), .a(\U1667/U1669/n2 ), .b(
        \U1667/U1669/nr ), .c(\U1667/U1669/nd ) );
    inv_2 \U1667/U1669/U3  ( .x(net193), .a(\U1667/U1669/n2 ) );
    buf_2 \U1650/U1653  ( .x(\U1650/latch ), .a(net172) );
    nor2_1 \U1650/U264/U5  ( .x(\U1650/nlocalcd ), .a(reset), .b(
        \U1650/localcd ) );
    nor2_1 \U1650/U1659_0_/U5  ( .x(\U1650/ncd[0] ), .a(\U1650/ol[0] ), .b(
        \U1650/oh[0] ) );
    nor2_1 \U1650/U1659_1_/U5  ( .x(\U1650/ncd[1] ), .a(\U1650/ol[1] ), .b(
        \U1650/oh[1] ) );
    nor2_1 \U1650/U1659_2_/U5  ( .x(\U1650/ncd[2] ), .a(\U1650/ol[2] ), .b(
        \U1650/oh[2] ) );
    nor2_1 \U1650/U1659_3_/U5  ( .x(\U1650/ncd[3] ), .a(\U1650/ol[3] ), .b(
        \U1650/oh[3] ) );
    nor2_1 \U1650/U1659_4_/U5  ( .x(\U1650/ncd[4] ), .a(\U1650/ol[4] ), .b(
        \U1650/oh[4] ) );
    nor2_1 \U1650/U1659_5_/U5  ( .x(\U1650/ncd[5] ), .a(\col_l[0] ), .b(
        \col_h[0] ) );
    nor2_1 \U1650/U1659_6_/U5  ( .x(\U1650/ncd[6] ), .a(\col_l[1] ), .b(
        \col_h[1] ) );
    nor2_1 \U1650/U1659_7_/U5  ( .x(\U1650/ncd[7] ), .a(\col_l[2] ), .b(
        \col_h[2] ) );
    nor2_1 \U1650/U3/U5  ( .x(\U1650/ctrlack_internal ), .a(\U1650/acb ), .b(
        \U1650/ba ) );
    buf_2 \U1650/U1665/U7  ( .x(\U1650/driveh ), .a(start_receiving) );
    buf_2 \U1650/U1666/U7  ( .x(\U1650/drivel ), .a(start_receiving) );
    ao23_1 \U1650/U1658_0_/U21/U1/U1  ( .x(\U1650/ol[0] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[0] ), .c(\U1650/drivel ), .d(cbl[0]), .e(n7) );
    ao23_1 \U1650/U1658_1_/U21/U1/U1  ( .x(\U1650/ol[1] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[1] ), .c(\U1650/drivel ), .d(cbl[1]), .e(n7) );
    ao23_1 \U1650/U1658_2_/U21/U1/U1  ( .x(\U1650/ol[2] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[2] ), .c(\U1650/drivel ), .d(cbl[2]), .e(n7) );
    ao23_1 \U1650/U1658_3_/U21/U1/U1  ( .x(\U1650/ol[3] ), .a(n9), .b(
        \U1650/ol[3] ), .c(\U1650/drivel ), .d(cbl[3]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1658_4_/U21/U1/U1  ( .x(\U1650/ol[4] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[4] ), .c(\U1650/drivel ), .d(cbl[4]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1658_5_/U21/U1/U1  ( .x(\col_l[0] ), .a(\U1650/drivel ), 
        .b(\col_l[0] ), .c(\U1650/drivel ), .d(cbl[5]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1658_6_/U21/U1/U1  ( .x(\col_l[1] ), .a(n9), .b(\col_l[1] ), 
        .c(\U1650/drivel ), .d(cbl[6]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1658_7_/U21/U1/U1  ( .x(\col_l[2] ), .a(n9), .b(\col_l[2] ), 
        .c(\U1650/drivel ), .d(cbl[7]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_0_/U21/U1/U1  ( .x(\U1650/oh[0] ), .a(\U1650/driveh ), 
        .b(\U1650/oh[0] ), .c(\U1650/driveh ), .d(cbh[0]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1651_1_/U21/U1/U1  ( .x(\U1650/oh[1] ), .a(\U1650/driveh ), 
        .b(\U1650/oh[1] ), .c(\U1650/driveh ), .d(cbh[1]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1651_2_/U21/U1/U1  ( .x(\U1650/oh[2] ), .a(\U1650/driveh ), 
        .b(\U1650/oh[2] ), .c(\U1650/driveh ), .d(cbh[2]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1651_3_/U21/U1/U1  ( .x(\U1650/oh[3] ), .a(n8), .b(
        \U1650/oh[3] ), .c(\U1650/driveh ), .d(cbh[3]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_4_/U21/U1/U1  ( .x(\U1650/oh[4] ), .a(n8), .b(
        \U1650/oh[4] ), .c(\U1650/driveh ), .d(cbh[4]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_5_/U21/U1/U1  ( .x(\col_h[0] ), .a(\U1650/driveh ), 
        .b(\col_h[0] ), .c(\U1650/driveh ), .d(cbh[5]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_6_/U21/U1/U1  ( .x(\col_h[1] ), .a(n8), .b(\col_h[1] ), 
        .c(\U1650/driveh ), .d(cbh[6]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_7_/U21/U1/U1  ( .x(\col_h[2] ), .a(\U1650/driveh ), 
        .b(\col_h[2] ), .c(\U1650/driveh ), .d(cbh[7]), .e(\U1650/latch ) );
    aoai211_1 \U1650/U4/U28/U1/U1  ( .x(\U1650/U4/U28/U1/clr ), .a(
        start_receiving), .b(\U1650/acb ), .c(\U1650/nlocalcd ), .d(net172) );
    nand3_1 \U1650/U4/U28/U1/U2  ( .x(\U1650/U4/U28/U1/set ), .a(
        \U1650/nlocalcd ), .b(start_receiving), .c(\U1650/acb ) );
    nand2_2 \U1650/U4/U28/U1/U3  ( .x(net172), .a(\U1650/U4/U28/U1/clr ), .b(
        \U1650/U4/U28/U1/set ) );
    oai21_1 \U1650/U1/U30/U1/U1  ( .x(\U1650/acb ), .a(\U1650/U1/Z ), .b(
        \U1650/ba ), .c(start_receiving) );
    inv_1 \U1650/U1/U30/U1/U2  ( .x(\U1650/U1/Z ), .a(\U1650/acb ) );
    ao222_1 \U1650/U5/U18/U1/U1  ( .x(\U1650/ba ), .a(\U1650/latch ), .b(n14), 
        .c(\U1650/latch ), .d(\U1650/ba ), .e(n14), .f(\U1650/ba ) );
    aoi222_1 \U1650/U1664/U28/U30/U1  ( .x(\U1650/U1664/x[3] ), .a(
        \U1650/ncd[7] ), .b(\U1650/ncd[6] ), .c(\U1650/ncd[7] ), .d(
        \U1650/U1664/U28/Z ), .e(\U1650/ncd[6] ), .f(\U1650/U1664/U28/Z ) );
    inv_1 \U1650/U1664/U28/U30/Uinv  ( .x(\U1650/U1664/U28/Z ), .a(
        \U1650/U1664/x[3] ) );
    aoi222_1 \U1650/U1664/U32/U30/U1  ( .x(\U1650/U1664/x[0] ), .a(
        \U1650/ncd[1] ), .b(\U1650/ncd[0] ), .c(\U1650/ncd[1] ), .d(
        \U1650/U1664/U32/Z ), .e(\U1650/ncd[0] ), .f(\U1650/U1664/U32/Z ) );
    inv_1 \U1650/U1664/U32/U30/Uinv  ( .x(\U1650/U1664/U32/Z ), .a(
        \U1650/U1664/x[0] ) );
    aoi222_1 \U1650/U1664/U29/U30/U1  ( .x(\U1650/U1664/x[2] ), .a(
        \U1650/ncd[5] ), .b(\U1650/ncd[4] ), .c(\U1650/ncd[5] ), .d(
        \U1650/U1664/U29/Z ), .e(\U1650/ncd[4] ), .f(\U1650/U1664/U29/Z ) );
    inv_1 \U1650/U1664/U29/U30/Uinv  ( .x(\U1650/U1664/U29/Z ), .a(
        \U1650/U1664/x[2] ) );
    aoi222_1 \U1650/U1664/U33/U30/U1  ( .x(\U1650/U1664/y[0] ), .a(
        \U1650/U1664/x[1] ), .b(\U1650/U1664/x[0] ), .c(\U1650/U1664/x[1] ), 
        .d(\U1650/U1664/U33/Z ), .e(\U1650/U1664/x[0] ), .f(
        \U1650/U1664/U33/Z ) );
    inv_1 \U1650/U1664/U33/U30/Uinv  ( .x(\U1650/U1664/U33/Z ), .a(
        \U1650/U1664/y[0] ) );
    aoi222_1 \U1650/U1664/U30/U30/U1  ( .x(\U1650/U1664/y[1] ), .a(
        \U1650/U1664/x[3] ), .b(\U1650/U1664/x[2] ), .c(\U1650/U1664/x[3] ), 
        .d(\U1650/U1664/U30/Z ), .e(\U1650/U1664/x[2] ), .f(
        \U1650/U1664/U30/Z ) );
    inv_1 \U1650/U1664/U30/U30/Uinv  ( .x(\U1650/U1664/U30/Z ), .a(
        \U1650/U1664/y[1] ) );
    aoi222_1 \U1650/U1664/U31/U30/U1  ( .x(\U1650/U1664/x[1] ), .a(
        \U1650/ncd[3] ), .b(\U1650/ncd[2] ), .c(\U1650/ncd[3] ), .d(
        \U1650/U1664/U31/Z ), .e(\U1650/ncd[2] ), .f(\U1650/U1664/U31/Z ) );
    inv_1 \U1650/U1664/U31/U30/Uinv  ( .x(\U1650/U1664/U31/Z ), .a(
        \U1650/U1664/x[1] ) );
    aoi222_1 \U1650/U1664/U37/U30/U1  ( .x(\U1650/localcd ), .a(
        \U1650/U1664/y[0] ), .b(\U1650/U1664/y[1] ), .c(\U1650/U1664/y[0] ), 
        .d(\U1650/U1664/U37/Z ), .e(\U1650/U1664/y[1] ), .f(
        \U1650/U1664/U37/Z ) );
    inv_1 \U1650/U1664/U37/U30/Uinv  ( .x(\U1650/U1664/U37/Z ), .a(
        \U1650/localcd ) );
    nor3_1 \U1650/U1669/Unr  ( .x(\U1650/U1669/nr ), .a(
        \U1650/ctrlack_internal ), .b(\U1650/drivel ), .c(\U1650/driveh ) );
    nand3_1 \U1650/U1669/Und  ( .x(\U1650/U1669/nd ), .a(
        \U1650/ctrlack_internal ), .b(\U1650/drivel ), .c(\U1650/driveh ) );
    oa21_1 \U1650/U1669/U1  ( .x(\U1650/U1669/n2 ), .a(\U1650/U1669/n2 ), .b(
        \U1650/U1669/nr ), .c(\U1650/U1669/nd ) );
    inv_2 \U1650/U1669/U3  ( .x(net139), .a(\U1650/U1669/n2 ) );
    buf_2 \U1666/U1653  ( .x(\U1666/latch ), .a(net169) );
    nor2_1 \U1666/U264/U5  ( .x(\U1666/nlocalcd ), .a(reset), .b(
        \U1666/localcd ) );
    nor2_1 \U1666/U1659_0_/U5  ( .x(\U1666/ncd[0] ), .a(rd[24]), .b(rd[56]) );
    nor2_1 \U1666/U1659_1_/U5  ( .x(\U1666/ncd[1] ), .a(rd[25]), .b(rd[57]) );
    nor2_1 \U1666/U1659_2_/U5  ( .x(\U1666/ncd[2] ), .a(rd[26]), .b(rd[58]) );
    nor2_1 \U1666/U1659_3_/U5  ( .x(\U1666/ncd[3] ), .a(rd[27]), .b(rd[59]) );
    nor2_1 \U1666/U1659_4_/U5  ( .x(\U1666/ncd[4] ), .a(rd[28]), .b(rd[60]) );
    nor2_1 \U1666/U1659_5_/U5  ( .x(\U1666/ncd[5] ), .a(rd[29]), .b(rd[61]) );
    nor2_1 \U1666/U1659_6_/U5  ( .x(\U1666/ncd[6] ), .a(rd[30]), .b(rd[62]) );
    nor2_1 \U1666/U1659_7_/U5  ( .x(\U1666/ncd[7] ), .a(rd[31]), .b(rd[63]) );
    nor2_1 \U1666/U3/U5  ( .x(\U1666/ctrlack_internal ), .a(\U1666/acb ), .b(
        \U1666/ba ) );
    buf_2 \U1666/U1665/U7  ( .x(\U1666/driveh ), .a(read) );
    buf_2 \U1666/U1666/U7  ( .x(\U1666/drivel ), .a(read) );
    ao23_1 \U1666/U1658_0_/U21/U1/U1  ( .x(rd[24]), .a(n6), .b(rd[24]), .c(
        \U1666/drivel ), .d(cbl[0]), .e(n5) );
    ao23_1 \U1666/U1658_1_/U21/U1/U1  ( .x(rd[25]), .a(n6), .b(rd[25]), .c(
        \U1666/driveh ), .d(cbl[1]), .e(n5) );
    ao23_1 \U1666/U1658_2_/U21/U1/U1  ( .x(rd[26]), .a(\U1666/driveh ), .b(rd
        [26]), .c(n6), .d(cbl[2]), .e(n5) );
    ao23_1 \U1666/U1658_3_/U21/U1/U1  ( .x(rd[27]), .a(n6), .b(rd[27]), .c(
        \U1666/driveh ), .d(cbl[3]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_4_/U21/U1/U1  ( .x(rd[28]), .a(\U1666/drivel ), .b(rd
        [28]), .c(n6), .d(cbl[4]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_5_/U21/U1/U1  ( .x(rd[29]), .a(\U1666/drivel ), .b(rd
        [29]), .c(n6), .d(cbl[5]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_6_/U21/U1/U1  ( .x(rd[30]), .a(\U1666/driveh ), .b(rd
        [30]), .c(\U1666/drivel ), .d(cbl[6]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_7_/U21/U1/U1  ( .x(rd[31]), .a(\U1666/driveh ), .b(rd
        [31]), .c(\U1666/driveh ), .d(cbl[7]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_0_/U21/U1/U1  ( .x(rd[56]), .a(\U1666/drivel ), .b(rd
        [56]), .c(n6), .d(cbh[0]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_1_/U21/U1/U1  ( .x(rd[57]), .a(\U1666/driveh ), .b(rd
        [57]), .c(\U1666/drivel ), .d(cbh[1]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_2_/U21/U1/U1  ( .x(rd[58]), .a(\U1666/drivel ), .b(rd
        [58]), .c(\U1666/drivel ), .d(cbh[2]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_3_/U21/U1/U1  ( .x(rd[59]), .a(\U1666/driveh ), .b(rd
        [59]), .c(\U1666/driveh ), .d(cbh[3]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_4_/U21/U1/U1  ( .x(rd[60]), .a(\U1666/drivel ), .b(rd
        [60]), .c(\U1666/driveh ), .d(cbh[4]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_5_/U21/U1/U1  ( .x(rd[61]), .a(\U1666/driveh ), .b(rd
        [61]), .c(n6), .d(cbh[5]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_6_/U21/U1/U1  ( .x(rd[62]), .a(n6), .b(rd[62]), .c(
        \U1666/drivel ), .d(cbh[6]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_7_/U21/U1/U1  ( .x(rd[63]), .a(n6), .b(rd[63]), .c(n6), 
        .d(cbh[7]), .e(\U1666/latch ) );
    aoai211_1 \U1666/U4/U28/U1/U1  ( .x(\U1666/U4/U28/U1/clr ), .a(read), .b(
        \U1666/acb ), .c(\U1666/nlocalcd ), .d(net169) );
    nand3_1 \U1666/U4/U28/U1/U2  ( .x(\U1666/U4/U28/U1/set ), .a(
        \U1666/nlocalcd ), .b(read), .c(\U1666/acb ) );
    nand2_2 \U1666/U4/U28/U1/U3  ( .x(net169), .a(\U1666/U4/U28/U1/clr ), .b(
        \U1666/U4/U28/U1/set ) );
    oai21_1 \U1666/U1/U30/U1/U1  ( .x(\U1666/acb ), .a(\U1666/U1/Z ), .b(
        \U1666/ba ), .c(read) );
    inv_1 \U1666/U1/U30/U1/U2  ( .x(\U1666/U1/Z ), .a(\U1666/acb ) );
    ao222_1 \U1666/U5/U18/U1/U1  ( .x(\U1666/ba ), .a(\U1666/latch ), .b(n14), 
        .c(\U1666/latch ), .d(\U1666/ba ), .e(n14), .f(\U1666/ba ) );
    aoi222_1 \U1666/U1664/U28/U30/U1  ( .x(\U1666/U1664/x[3] ), .a(
        \U1666/ncd[7] ), .b(\U1666/ncd[6] ), .c(\U1666/ncd[7] ), .d(
        \U1666/U1664/U28/Z ), .e(\U1666/ncd[6] ), .f(\U1666/U1664/U28/Z ) );
    inv_1 \U1666/U1664/U28/U30/Uinv  ( .x(\U1666/U1664/U28/Z ), .a(
        \U1666/U1664/x[3] ) );
    aoi222_1 \U1666/U1664/U32/U30/U1  ( .x(\U1666/U1664/x[0] ), .a(
        \U1666/ncd[1] ), .b(\U1666/ncd[0] ), .c(\U1666/ncd[1] ), .d(
        \U1666/U1664/U32/Z ), .e(\U1666/ncd[0] ), .f(\U1666/U1664/U32/Z ) );
    inv_1 \U1666/U1664/U32/U30/Uinv  ( .x(\U1666/U1664/U32/Z ), .a(
        \U1666/U1664/x[0] ) );
    aoi222_1 \U1666/U1664/U29/U30/U1  ( .x(\U1666/U1664/x[2] ), .a(
        \U1666/ncd[5] ), .b(\U1666/ncd[4] ), .c(\U1666/ncd[5] ), .d(
        \U1666/U1664/U29/Z ), .e(\U1666/ncd[4] ), .f(\U1666/U1664/U29/Z ) );
    inv_1 \U1666/U1664/U29/U30/Uinv  ( .x(\U1666/U1664/U29/Z ), .a(
        \U1666/U1664/x[2] ) );
    aoi222_1 \U1666/U1664/U33/U30/U1  ( .x(\U1666/U1664/y[0] ), .a(
        \U1666/U1664/x[1] ), .b(\U1666/U1664/x[0] ), .c(\U1666/U1664/x[1] ), 
        .d(\U1666/U1664/U33/Z ), .e(\U1666/U1664/x[0] ), .f(
        \U1666/U1664/U33/Z ) );
    inv_1 \U1666/U1664/U33/U30/Uinv  ( .x(\U1666/U1664/U33/Z ), .a(
        \U1666/U1664/y[0] ) );
    aoi222_1 \U1666/U1664/U30/U30/U1  ( .x(\U1666/U1664/y[1] ), .a(
        \U1666/U1664/x[3] ), .b(\U1666/U1664/x[2] ), .c(\U1666/U1664/x[3] ), 
        .d(\U1666/U1664/U30/Z ), .e(\U1666/U1664/x[2] ), .f(
        \U1666/U1664/U30/Z ) );
    inv_1 \U1666/U1664/U30/U30/Uinv  ( .x(\U1666/U1664/U30/Z ), .a(
        \U1666/U1664/y[1] ) );
    aoi222_1 \U1666/U1664/U31/U30/U1  ( .x(\U1666/U1664/x[1] ), .a(
        \U1666/ncd[3] ), .b(\U1666/ncd[2] ), .c(\U1666/ncd[3] ), .d(
        \U1666/U1664/U31/Z ), .e(\U1666/ncd[2] ), .f(\U1666/U1664/U31/Z ) );
    inv_1 \U1666/U1664/U31/U30/Uinv  ( .x(\U1666/U1664/U31/Z ), .a(
        \U1666/U1664/x[1] ) );
    aoi222_1 \U1666/U1664/U37/U30/U1  ( .x(\U1666/localcd ), .a(
        \U1666/U1664/y[0] ), .b(\U1666/U1664/y[1] ), .c(\U1666/U1664/y[0] ), 
        .d(\U1666/U1664/U37/Z ), .e(\U1666/U1664/y[1] ), .f(
        \U1666/U1664/U37/Z ) );
    inv_1 \U1666/U1664/U37/U30/Uinv  ( .x(\U1666/U1664/U37/Z ), .a(
        \U1666/localcd ) );
    nor3_1 \U1666/U1669/Unr  ( .x(\U1666/U1669/nr ), .a(
        \U1666/ctrlack_internal ), .b(n6), .c(\U1666/drivel ) );
    nand3_1 \U1666/U1669/Und  ( .x(\U1666/U1669/nd ), .a(
        \U1666/ctrlack_internal ), .b(\U1666/driveh ), .c(\U1666/drivel ) );
    oa21_1 \U1666/U1669/U1  ( .x(\U1666/U1669/n2 ), .a(\U1666/U1669/n2 ), .b(
        \U1666/U1669/nr ), .c(\U1666/U1669/nd ) );
    inv_2 \U1666/U1669/U3  ( .x(net94), .a(\U1666/U1669/n2 ) );
    buf_2 \I1/U1653  ( .x(\I1/latch ), .a(net166) );
    nor2_1 \I1/U264/U5  ( .x(\I1/nlocalcd ), .a(reset), .b(\I1/localcd ) );
    nor2_1 \I1/U1659_0_/U5  ( .x(\I1/ncd[0] ), .a(rd[8]), .b(rd[40]) );
    nor2_1 \I1/U1659_1_/U5  ( .x(\I1/ncd[1] ), .a(rd[9]), .b(rd[41]) );
    nor2_1 \I1/U1659_2_/U5  ( .x(\I1/ncd[2] ), .a(rd[10]), .b(rd[42]) );
    nor2_1 \I1/U1659_3_/U5  ( .x(\I1/ncd[3] ), .a(rd[11]), .b(rd[43]) );
    nor2_1 \I1/U1659_4_/U5  ( .x(\I1/ncd[4] ), .a(rd[12]), .b(rd[44]) );
    nor2_1 \I1/U1659_5_/U5  ( .x(\I1/ncd[5] ), .a(rd[13]), .b(rd[45]) );
    nor2_1 \I1/U1659_6_/U5  ( .x(\I1/ncd[6] ), .a(rd[14]), .b(rd[46]) );
    nor2_1 \I1/U1659_7_/U5  ( .x(\I1/ncd[7] ), .a(rd[15]), .b(rd[47]) );
    nor2_1 \I1/U3/U5  ( .x(\I1/ctrlack_internal ), .a(\I1/acb ), .b(\I1/ba )
         );
    buf_2 \I1/U1665/U7  ( .x(\I1/driveh ), .a(net103) );
    buf_2 \I1/U1666/U7  ( .x(\I1/drivel ), .a(net103) );
    ao23_1 \I1/U1658_0_/U21/U1/U1  ( .x(rd[8]), .a(n4), .b(rd[8]), .c(
        \I1/drivel ), .d(cbl[0]), .e(n3) );
    ao23_1 \I1/U1658_1_/U21/U1/U1  ( .x(rd[9]), .a(n4), .b(rd[9]), .c(
        \I1/driveh ), .d(cbl[1]), .e(n3) );
    ao23_1 \I1/U1658_2_/U21/U1/U1  ( .x(rd[10]), .a(\I1/driveh ), .b(rd[10]), 
        .c(n4), .d(cbl[2]), .e(n3) );
    ao23_1 \I1/U1658_3_/U21/U1/U1  ( .x(rd[11]), .a(n4), .b(rd[11]), .c(
        \I1/driveh ), .d(cbl[3]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_4_/U21/U1/U1  ( .x(rd[12]), .a(\I1/drivel ), .b(rd[12]), 
        .c(n4), .d(cbl[4]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_5_/U21/U1/U1  ( .x(rd[13]), .a(\I1/drivel ), .b(rd[13]), 
        .c(n4), .d(cbl[5]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_6_/U21/U1/U1  ( .x(rd[14]), .a(\I1/driveh ), .b(rd[14]), 
        .c(\I1/drivel ), .d(cbl[6]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_7_/U21/U1/U1  ( .x(rd[15]), .a(\I1/driveh ), .b(rd[15]), 
        .c(\I1/driveh ), .d(cbl[7]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_0_/U21/U1/U1  ( .x(rd[40]), .a(\I1/drivel ), .b(rd[40]), 
        .c(n4), .d(cbh[0]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_1_/U21/U1/U1  ( .x(rd[41]), .a(\I1/driveh ), .b(rd[41]), 
        .c(\I1/drivel ), .d(cbh[1]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_2_/U21/U1/U1  ( .x(rd[42]), .a(\I1/drivel ), .b(rd[42]), 
        .c(\I1/drivel ), .d(cbh[2]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_3_/U21/U1/U1  ( .x(rd[43]), .a(\I1/driveh ), .b(rd[43]), 
        .c(\I1/driveh ), .d(cbh[3]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_4_/U21/U1/U1  ( .x(rd[44]), .a(\I1/drivel ), .b(rd[44]), 
        .c(\I1/driveh ), .d(cbh[4]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_5_/U21/U1/U1  ( .x(rd[45]), .a(\I1/driveh ), .b(rd[45]), 
        .c(n4), .d(cbh[5]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_6_/U21/U1/U1  ( .x(rd[46]), .a(n4), .b(rd[46]), .c(
        \I1/drivel ), .d(cbh[6]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_7_/U21/U1/U1  ( .x(rd[47]), .a(n4), .b(rd[47]), .c(n4), 
        .d(cbh[7]), .e(\I1/latch ) );
    aoai211_1 \I1/U4/U28/U1/U1  ( .x(\I1/U4/U28/U1/clr ), .a(net103), .b(
        \I1/acb ), .c(\I1/nlocalcd ), .d(net166) );
    nand3_1 \I1/U4/U28/U1/U2  ( .x(\I1/U4/U28/U1/set ), .a(\I1/nlocalcd ), .b(
        net103), .c(\I1/acb ) );
    nand2_2 \I1/U4/U28/U1/U3  ( .x(net166), .a(\I1/U4/U28/U1/clr ), .b(
        \I1/U4/U28/U1/set ) );
    oai21_1 \I1/U1/U30/U1/U1  ( .x(\I1/acb ), .a(\I1/U1/Z ), .b(\I1/ba ), .c(
        net103) );
    inv_1 \I1/U1/U30/U1/U2  ( .x(\I1/U1/Z ), .a(\I1/acb ) );
    ao222_1 \I1/U5/U18/U1/U1  ( .x(\I1/ba ), .a(\I1/latch ), .b(n14), .c(
        \I1/latch ), .d(\I1/ba ), .e(n14), .f(\I1/ba ) );
    aoi222_1 \I1/U1664/U28/U30/U1  ( .x(\I1/U1664/x[3] ), .a(\I1/ncd[7] ), .b(
        \I1/ncd[6] ), .c(\I1/ncd[7] ), .d(\I1/U1664/U28/Z ), .e(\I1/ncd[6] ), 
        .f(\I1/U1664/U28/Z ) );
    inv_1 \I1/U1664/U28/U30/Uinv  ( .x(\I1/U1664/U28/Z ), .a(\I1/U1664/x[3] )
         );
    aoi222_1 \I1/U1664/U32/U30/U1  ( .x(\I1/U1664/x[0] ), .a(\I1/ncd[1] ), .b(
        \I1/ncd[0] ), .c(\I1/ncd[1] ), .d(\I1/U1664/U32/Z ), .e(\I1/ncd[0] ), 
        .f(\I1/U1664/U32/Z ) );
    inv_1 \I1/U1664/U32/U30/Uinv  ( .x(\I1/U1664/U32/Z ), .a(\I1/U1664/x[0] )
         );
    aoi222_1 \I1/U1664/U29/U30/U1  ( .x(\I1/U1664/x[2] ), .a(\I1/ncd[5] ), .b(
        \I1/ncd[4] ), .c(\I1/ncd[5] ), .d(\I1/U1664/U29/Z ), .e(\I1/ncd[4] ), 
        .f(\I1/U1664/U29/Z ) );
    inv_1 \I1/U1664/U29/U30/Uinv  ( .x(\I1/U1664/U29/Z ), .a(\I1/U1664/x[2] )
         );
    aoi222_1 \I1/U1664/U33/U30/U1  ( .x(\I1/U1664/y[0] ), .a(\I1/U1664/x[1] ), 
        .b(\I1/U1664/x[0] ), .c(\I1/U1664/x[1] ), .d(\I1/U1664/U33/Z ), .e(
        \I1/U1664/x[0] ), .f(\I1/U1664/U33/Z ) );
    inv_1 \I1/U1664/U33/U30/Uinv  ( .x(\I1/U1664/U33/Z ), .a(\I1/U1664/y[0] )
         );
    aoi222_1 \I1/U1664/U30/U30/U1  ( .x(\I1/U1664/y[1] ), .a(\I1/U1664/x[3] ), 
        .b(\I1/U1664/x[2] ), .c(\I1/U1664/x[3] ), .d(\I1/U1664/U30/Z ), .e(
        \I1/U1664/x[2] ), .f(\I1/U1664/U30/Z ) );
    inv_1 \I1/U1664/U30/U30/Uinv  ( .x(\I1/U1664/U30/Z ), .a(\I1/U1664/y[1] )
         );
    aoi222_1 \I1/U1664/U31/U30/U1  ( .x(\I1/U1664/x[1] ), .a(\I1/ncd[3] ), .b(
        \I1/ncd[2] ), .c(\I1/ncd[3] ), .d(\I1/U1664/U31/Z ), .e(\I1/ncd[2] ), 
        .f(\I1/U1664/U31/Z ) );
    inv_1 \I1/U1664/U31/U30/Uinv  ( .x(\I1/U1664/U31/Z ), .a(\I1/U1664/x[1] )
         );
    aoi222_1 \I1/U1664/U37/U30/U1  ( .x(\I1/localcd ), .a(\I1/U1664/y[0] ), 
        .b(\I1/U1664/y[1] ), .c(\I1/U1664/y[0] ), .d(\I1/U1664/U37/Z ), .e(
        \I1/U1664/y[1] ), .f(\I1/U1664/U37/Z ) );
    inv_1 \I1/U1664/U37/U30/Uinv  ( .x(\I1/U1664/U37/Z ), .a(\I1/localcd ) );
    nor3_1 \I1/U1669/Unr  ( .x(\I1/U1669/nr ), .a(\I1/ctrlack_internal ), .b(
        n4), .c(\I1/drivel ) );
    nand3_1 \I1/U1669/Und  ( .x(\I1/U1669/nd ), .a(\I1/ctrlack_internal ), .b(
        \I1/driveh ), .c(\I1/drivel ) );
    oa21_1 \I1/U1669/U1  ( .x(\I1/U1669/n2 ), .a(\I1/U1669/n2 ), .b(
        \I1/U1669/nr ), .c(\I1/U1669/nd ) );
    inv_2 \I1/U1669/U3  ( .x(read_lhw), .a(\I1/U1669/n2 ) );
    buf_2 \I2/U1653  ( .x(\I2/latch ), .a(net170) );
    nor2_1 \I2/U264/U5  ( .x(\I2/nlocalcd ), .a(reset), .b(\I2/localcd ) );
    nor2_1 \I2/U1659_0_/U5  ( .x(\I2/ncd[0] ), .a(rd[16]), .b(rd[48]) );
    nor2_1 \I2/U1659_1_/U5  ( .x(\I2/ncd[1] ), .a(rd[17]), .b(rd[49]) );
    nor2_1 \I2/U1659_2_/U5  ( .x(\I2/ncd[2] ), .a(rd[18]), .b(rd[50]) );
    nor2_1 \I2/U1659_3_/U5  ( .x(\I2/ncd[3] ), .a(rd[19]), .b(rd[51]) );
    nor2_1 \I2/U1659_4_/U5  ( .x(\I2/ncd[4] ), .a(rd[20]), .b(rd[52]) );
    nor2_1 \I2/U1659_5_/U5  ( .x(\I2/ncd[5] ), .a(rd[21]), .b(rd[53]) );
    nor2_1 \I2/U1659_6_/U5  ( .x(\I2/ncd[6] ), .a(rd[22]), .b(rd[54]) );
    nor2_1 \I2/U1659_7_/U5  ( .x(\I2/ncd[7] ), .a(rd[23]), .b(rd[55]) );
    nor2_1 \I2/U3/U5  ( .x(\I2/ctrlack_internal ), .a(\I2/acb ), .b(\I2/ba )
         );
    buf_2 \I2/U1665/U7  ( .x(\I2/driveh ), .a(net94) );
    buf_2 \I2/U1666/U7  ( .x(\I2/drivel ), .a(net94) );
    ao23_1 \I2/U1658_0_/U21/U1/U1  ( .x(rd[16]), .a(n2), .b(rd[16]), .c(
        \I2/drivel ), .d(cbl[0]), .e(n1) );
    ao23_1 \I2/U1658_1_/U21/U1/U1  ( .x(rd[17]), .a(n2), .b(rd[17]), .c(
        \I2/driveh ), .d(cbl[1]), .e(n1) );
    ao23_1 \I2/U1658_2_/U21/U1/U1  ( .x(rd[18]), .a(\I2/driveh ), .b(rd[18]), 
        .c(n2), .d(cbl[2]), .e(n1) );
    ao23_1 \I2/U1658_3_/U21/U1/U1  ( .x(rd[19]), .a(n2), .b(rd[19]), .c(
        \I2/driveh ), .d(cbl[3]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_4_/U21/U1/U1  ( .x(rd[20]), .a(\I2/drivel ), .b(rd[20]), 
        .c(n2), .d(cbl[4]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_5_/U21/U1/U1  ( .x(rd[21]), .a(\I2/drivel ), .b(rd[21]), 
        .c(n2), .d(cbl[5]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_6_/U21/U1/U1  ( .x(rd[22]), .a(\I2/driveh ), .b(rd[22]), 
        .c(\I2/drivel ), .d(cbl[6]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_7_/U21/U1/U1  ( .x(rd[23]), .a(\I2/driveh ), .b(rd[23]), 
        .c(\I2/driveh ), .d(cbl[7]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_0_/U21/U1/U1  ( .x(rd[48]), .a(\I2/drivel ), .b(rd[48]), 
        .c(n2), .d(cbh[0]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_1_/U21/U1/U1  ( .x(rd[49]), .a(\I2/driveh ), .b(rd[49]), 
        .c(\I2/drivel ), .d(cbh[1]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_2_/U21/U1/U1  ( .x(rd[50]), .a(\I2/drivel ), .b(rd[50]), 
        .c(\I2/drivel ), .d(cbh[2]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_3_/U21/U1/U1  ( .x(rd[51]), .a(\I2/driveh ), .b(rd[51]), 
        .c(\I2/driveh ), .d(cbh[3]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_4_/U21/U1/U1  ( .x(rd[52]), .a(\I2/drivel ), .b(rd[52]), 
        .c(\I2/driveh ), .d(cbh[4]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_5_/U21/U1/U1  ( .x(rd[53]), .a(\I2/driveh ), .b(rd[53]), 
        .c(n2), .d(cbh[5]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_6_/U21/U1/U1  ( .x(rd[54]), .a(n2), .b(rd[54]), .c(
        \I2/drivel ), .d(cbh[6]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_7_/U21/U1/U1  ( .x(rd[55]), .a(n2), .b(rd[55]), .c(n2), 
        .d(cbh[7]), .e(\I2/latch ) );
    aoai211_1 \I2/U4/U28/U1/U1  ( .x(\I2/U4/U28/U1/clr ), .a(net94), .b(
        \I2/acb ), .c(\I2/nlocalcd ), .d(net170) );
    nand3_1 \I2/U4/U28/U1/U2  ( .x(\I2/U4/U28/U1/set ), .a(\I2/nlocalcd ), .b(
        net94), .c(\I2/acb ) );
    nand2_2 \I2/U4/U28/U1/U3  ( .x(net170), .a(\I2/U4/U28/U1/clr ), .b(
        \I2/U4/U28/U1/set ) );
    oai21_1 \I2/U1/U30/U1/U1  ( .x(\I2/acb ), .a(\I2/U1/Z ), .b(\I2/ba ), .c(
        net94) );
    inv_1 \I2/U1/U30/U1/U2  ( .x(\I2/U1/Z ), .a(\I2/acb ) );
    ao222_1 \I2/U5/U18/U1/U1  ( .x(\I2/ba ), .a(\I2/latch ), .b(n14), .c(
        \I2/latch ), .d(\I2/ba ), .e(n14), .f(\I2/ba ) );
    aoi222_1 \I2/U1664/U28/U30/U1  ( .x(\I2/U1664/x[3] ), .a(\I2/ncd[7] ), .b(
        \I2/ncd[6] ), .c(\I2/ncd[7] ), .d(\I2/U1664/U28/Z ), .e(\I2/ncd[6] ), 
        .f(\I2/U1664/U28/Z ) );
    inv_1 \I2/U1664/U28/U30/Uinv  ( .x(\I2/U1664/U28/Z ), .a(\I2/U1664/x[3] )
         );
    aoi222_1 \I2/U1664/U32/U30/U1  ( .x(\I2/U1664/x[0] ), .a(\I2/ncd[1] ), .b(
        \I2/ncd[0] ), .c(\I2/ncd[1] ), .d(\I2/U1664/U32/Z ), .e(\I2/ncd[0] ), 
        .f(\I2/U1664/U32/Z ) );
    inv_1 \I2/U1664/U32/U30/Uinv  ( .x(\I2/U1664/U32/Z ), .a(\I2/U1664/x[0] )
         );
    aoi222_1 \I2/U1664/U29/U30/U1  ( .x(\I2/U1664/x[2] ), .a(\I2/ncd[5] ), .b(
        \I2/ncd[4] ), .c(\I2/ncd[5] ), .d(\I2/U1664/U29/Z ), .e(\I2/ncd[4] ), 
        .f(\I2/U1664/U29/Z ) );
    inv_1 \I2/U1664/U29/U30/Uinv  ( .x(\I2/U1664/U29/Z ), .a(\I2/U1664/x[2] )
         );
    aoi222_1 \I2/U1664/U33/U30/U1  ( .x(\I2/U1664/y[0] ), .a(\I2/U1664/x[1] ), 
        .b(\I2/U1664/x[0] ), .c(\I2/U1664/x[1] ), .d(\I2/U1664/U33/Z ), .e(
        \I2/U1664/x[0] ), .f(\I2/U1664/U33/Z ) );
    inv_1 \I2/U1664/U33/U30/Uinv  ( .x(\I2/U1664/U33/Z ), .a(\I2/U1664/y[0] )
         );
    aoi222_1 \I2/U1664/U30/U30/U1  ( .x(\I2/U1664/y[1] ), .a(\I2/U1664/x[3] ), 
        .b(\I2/U1664/x[2] ), .c(\I2/U1664/x[3] ), .d(\I2/U1664/U30/Z ), .e(
        \I2/U1664/x[2] ), .f(\I2/U1664/U30/Z ) );
    inv_1 \I2/U1664/U30/U30/Uinv  ( .x(\I2/U1664/U30/Z ), .a(\I2/U1664/y[1] )
         );
    aoi222_1 \I2/U1664/U31/U30/U1  ( .x(\I2/U1664/x[1] ), .a(\I2/ncd[3] ), .b(
        \I2/ncd[2] ), .c(\I2/ncd[3] ), .d(\I2/U1664/U31/Z ), .e(\I2/ncd[2] ), 
        .f(\I2/U1664/U31/Z ) );
    inv_1 \I2/U1664/U31/U30/Uinv  ( .x(\I2/U1664/U31/Z ), .a(\I2/U1664/x[1] )
         );
    aoi222_1 \I2/U1664/U37/U30/U1  ( .x(\I2/localcd ), .a(\I2/U1664/y[0] ), 
        .b(\I2/U1664/y[1] ), .c(\I2/U1664/y[0] ), .d(\I2/U1664/U37/Z ), .e(
        \I2/U1664/y[1] ), .f(\I2/U1664/U37/Z ) );
    inv_1 \I2/U1664/U37/U30/Uinv  ( .x(\I2/U1664/U37/Z ), .a(\I2/localcd ) );
    nor3_1 \I2/U1669/Unr  ( .x(\I2/U1669/nr ), .a(\I2/ctrlack_internal ), .b(
        n2), .c(\I2/drivel ) );
    nand3_1 \I2/U1669/Und  ( .x(\I2/U1669/nd ), .a(\I2/ctrlack_internal ), .b(
        \I2/driveh ), .c(\I2/drivel ) );
    oa21_1 \I2/U1669/U1  ( .x(\I2/U1669/n2 ), .a(\I2/U1669/n2 ), .b(
        \I2/U1669/nr ), .c(\I2/U1669/nd ) );
    inv_2 \I2/U1669/U3  ( .x(net103), .a(\I2/U1669/n2 ) );
    buf_1 U1 ( .x(n1), .a(\I2/latch ) );
    buf_2 U2 ( .x(n2), .a(net94) );
    buf_1 U3 ( .x(n3), .a(\I1/latch ) );
    buf_2 U4 ( .x(n4), .a(net103) );
    buf_1 U5 ( .x(n5), .a(\U1666/latch ) );
    buf_2 U6 ( .x(n6), .a(read) );
    buf_1 U7 ( .x(n7), .a(\U1650/latch ) );
    buf_1 U8 ( .x(n8), .a(\U1650/driveh ) );
    buf_1 U9 ( .x(n9), .a(\U1650/drivel ) );
    buf_1 U10 ( .x(n10), .a(\U1667/latch ) );
    buf_2 U11 ( .x(n11), .a(read_lhw) );
    buf_1 U12 ( .x(n12), .a(\I6/latch ) );
    buf_2 U13 ( .x(n13), .a(net139) );
    buf_3 U14 ( .x(n14), .a(bpullcd) );
    buf_3 U15 ( .x(err[1]), .a(n17) );
    buf_3 U16 ( .x(err[0]), .a(n18) );
endmodule


module chain_fr2dr_byte_4 ( nia, oh, ol, i, nReset, noa );
output [7:0] oh;
output [7:0] ol;
input  [4:0] i;
input  nReset, noa;
output nia;
    wire eop, net135, nca, nbReset, ncla, \c[3] , \c[2] , \c[1] , \c[0] , 
        \cl[3] , \cl[2] , \cl[1] , \cl[0] , asel, bsel, asela, bsela, csel, 
        dsel, csela, dsela, esel, fsel, esela, fsela, naa, nda, \a[3] , \a[2] , 
        \a[1] , \a[0] , \d[3] , \d[2] , \d[1] , \d[0] , nba, nea, nfa, \b[3] , 
        \b[2] , \b[1] , \b[0] , \f[3] , \f[2] , \f[1] , \f[0] , \e[3] , \e[2] , 
        \e[1] , \e[0] , \U891/nack , \U891/acka , \U891/naack[0] , 
        \U891/naack[1] , \U891/iay , \U891/ackb , \U891/reset , \U891/neopack , 
        \U891/U1128/nb , \U891/U1128/na , \U891/U1118_0_/nr , 
        \U891/U1118_0_/nd , \U891/U1118_0_/n2 , \U891/U1118_1_/nr , 
        \U891/U1118_1_/nd , \U891/U1118_1_/n2 , \U891/U1118_2_/nr , 
        \U891/U1118_2_/nd , \U891/U1118_2_/n2 , \U891/U1118_3_/nr , 
        \U891/U1118_3_/nd , \U891/U1118_3_/n2 , \U891/U1117_0_/nr , 
        \U891/U1117_0_/nd , \U891/U1117_0_/n2 , \U891/U1117_1_/nr , 
        \U891/U1117_1_/nd , \U891/U1117_1_/n2 , \U891/U1117_2_/nr , 
        \U891/U1117_2_/nd , \U891/U1117_2_/n2 , \U891/U1117_3_/nr , 
        \U891/U1117_3_/nd , \U891/U1117_3_/n2 , \U886/nack , \U886/acka , 
        \U886/ackb , \U886/reset , \U886/U1128/nb , \U886/U1128/na , 
        \U886/U1127/n5 , \U886/U1127/n1 , \U886/U1127/n2 , \U886/U1127/n3 , 
        \U886/U1127/n4 , \U886/U1118_0_/nr , \U886/U1118_0_/nd , 
        \U886/U1118_0_/n2 , \U886/U1118_1_/nr , \U886/U1118_1_/nd , 
        \U886/U1118_1_/n2 , \U886/U1118_2_/nr , \U886/U1118_2_/nd , 
        \U886/U1118_2_/n2 , \U886/U1118_3_/nr , \U886/U1118_3_/nd , 
        \U886/U1118_3_/n2 , \U886/U1117_0_/nr , \U886/U1117_0_/nd , 
        \U886/U1117_0_/n2 , \U886/U1117_1_/nr , \U886/U1117_1_/nd , 
        \U886/U1117_1_/n2 , \U886/U1117_2_/nr , \U886/U1117_2_/nd , 
        \U886/U1117_2_/n2 , \U886/U1117_3_/nr , \U886/U1117_3_/nd , 
        \U886/U1117_3_/n2 , \U884/nack , \U884/acka , \U884/ackb , 
        \U884/reset , \U884/U1128/nb , \U884/U1128/na , \U884/U1127/n5 , 
        \U884/U1127/n1 , \U884/U1127/n2 , \U884/U1127/n3 , \U884/U1127/n4 , 
        \U884/U1118_0_/nr , \U884/U1118_0_/nd , \U884/U1118_0_/n2 , 
        \U884/U1118_1_/nr , \U884/U1118_1_/nd , \U884/U1118_1_/n2 , 
        \U884/U1118_2_/nr , \U884/U1118_2_/nd , \U884/U1118_2_/n2 , 
        \U884/U1118_3_/nr , \U884/U1118_3_/nd , \U884/U1118_3_/n2 , 
        \U884/U1117_0_/nr , \U884/U1117_0_/nd , \U884/U1117_0_/n2 , 
        \U884/U1117_1_/nr , \U884/U1117_1_/nd , \U884/U1117_1_/n2 , 
        \U884/U1117_2_/nr , \U884/U1117_2_/nd , \U884/U1117_2_/n2 , 
        \U884/U1117_3_/nr , \U884/U1117_3_/nd , \U884/U1117_3_/n2 , 
        \U888/naack , \U888/r , \U888/s , \U888/nback , \U888/reset , 
        \U887/naack , \U887/r , \U887/s , \U887/nback , \U887/reset , 
        \U885/naack , \U885/r , \U885/s , \U885/nback , \U885/reset , \U877/x , 
        \U877/y , \U877/reset , \U877/U590/U25/U1/clr , \U877/U590/U25/U1/ob , 
        \U877/U589/U25/U1/clr , \U877/U589/U25/U1/ob , \U877/U588/U25/U1/clr , 
        \U877/U588/U25/U1/ob , \U877/U591/U25/U1/clr , \U877/U591/U25/U1/ob , 
        \U876/x , \U876/y , \U876/reset , \U876/U590/U25/U1/clr , 
        \U876/U590/U25/U1/ob , \U876/U589/U25/U1/clr , \U876/U589/U25/U1/ob , 
        \U876/U588/U25/U1/clr , \U876/U588/U25/U1/ob , \U876/U591/U25/U1/clr , 
        \U876/U591/U25/U1/ob , \U2/x , \U2/y , \U2/reset , 
        \U2/U590/U25/U1/clr , \U2/U590/U25/U1/ob , \U2/U589/U25/U1/clr , 
        \U2/U589/U25/U1/ob , \U2/U588/U25/U1/clr , \U2/U588/U25/U1/ob , 
        \U2/U591/U25/U1/clr , \U2/U591/U25/U1/ob , \U1/x , \U1/y , \U1/reset , 
        \U1/U590/U25/U1/clr , \U1/U590/U25/U1/ob , \U1/U589/U25/U1/clr , 
        \U1/U589/U25/U1/ob , \U1/U588/U25/U1/clr , \U1/U588/U25/U1/ob , 
        \U1/U591/U25/U1/clr , \U1/U591/U25/U1/ob , \U881/nack[1] , 
        \U881/nack[0] , n1;
    buf_2 U897 ( .x(nbReset), .a(nReset) );
    and4_1 \U894/U12  ( .x(eop), .a(ncla), .b(csela), .c(asela), .d(i[4]) );
    inv_1 \U891/U1126/U3  ( .x(\U891/reset ), .a(nbReset) );
    inv_1 \U891/U1139/U3  ( .x(\U891/neopack ), .a(eop) );
    nand3_1 \U891/U1131/U9  ( .x(\U891/iay ), .a(\U891/neopack ), .b(
        \U891/naack[0] ), .c(\U891/naack[1] ) );
    nor3_1 \U891/U1128/U27  ( .x(\U891/U1128/nb ), .a(\U891/reset ), .b(\b[3] 
        ), .c(\b[2] ) );
    nor2_1 \U891/U1128/U26  ( .x(\U891/U1128/na ), .a(\b[1] ), .b(\b[0] ) );
    nand2_2 \U891/U1128/U29  ( .x(\U891/ackb ), .a(\U891/U1128/nb ), .b(
        \U891/U1128/na ) );
    nor2_1 \U891/U1133/U5  ( .x(\U891/naack[0] ), .a(\a[3] ), .b(\a[2] ) );
    nor2_1 \U891/U1108/U5  ( .x(\U891/nack ), .a(\U891/acka ), .b(\U891/ackb )
         );
    nor2_1 \U891/U1134/U5  ( .x(\U891/naack[1] ), .a(\a[1] ), .b(\a[0] ) );
    nor2_2 \U891/U914/U6  ( .x(nia), .a(\U891/iay ), .b(\U891/ackb ) );
    nand2_1 \U891/U1130/U5  ( .x(\U891/acka ), .a(\U891/naack[0] ), .b(
        \U891/naack[1] ) );
    ao222_4 \U891/U1121/U1/U1  ( .x(bsela), .a(\U891/nack ), .b(bsel), .c(
        \U891/nack ), .d(bsela), .e(bsel), .f(bsela) );
    ao222_4 \U891/U1120/U1/U1  ( .x(asela), .a(asel), .b(\U891/nack ), .c(asel
        ), .d(asela), .e(\U891/nack ), .f(asela) );
    nor3_1 \U891/U1118_0_/Unr  ( .x(\U891/U1118_0_/nr ), .a(i[0]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_0_/Und  ( .x(\U891/U1118_0_/nd ), .a(i[0]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_0_/U1  ( .x(\U891/U1118_0_/n2 ), .a(\U891/U1118_0_/n2 ), 
        .b(\U891/U1118_0_/nr ), .c(\U891/U1118_0_/nd ) );
    inv_2 \U891/U1118_0_/U3  ( .x(\a[0] ), .a(\U891/U1118_0_/n2 ) );
    nor3_1 \U891/U1118_1_/Unr  ( .x(\U891/U1118_1_/nr ), .a(i[1]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_1_/Und  ( .x(\U891/U1118_1_/nd ), .a(i[1]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_1_/U1  ( .x(\U891/U1118_1_/n2 ), .a(\U891/U1118_1_/n2 ), 
        .b(\U891/U1118_1_/nr ), .c(\U891/U1118_1_/nd ) );
    inv_2 \U891/U1118_1_/U3  ( .x(\a[1] ), .a(\U891/U1118_1_/n2 ) );
    nor3_1 \U891/U1118_2_/Unr  ( .x(\U891/U1118_2_/nr ), .a(i[2]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_2_/Und  ( .x(\U891/U1118_2_/nd ), .a(i[2]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_2_/U1  ( .x(\U891/U1118_2_/n2 ), .a(\U891/U1118_2_/n2 ), 
        .b(\U891/U1118_2_/nr ), .c(\U891/U1118_2_/nd ) );
    inv_2 \U891/U1118_2_/U3  ( .x(\a[2] ), .a(\U891/U1118_2_/n2 ) );
    nor3_1 \U891/U1118_3_/Unr  ( .x(\U891/U1118_3_/nr ), .a(i[3]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_3_/Und  ( .x(\U891/U1118_3_/nd ), .a(i[3]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_3_/U1  ( .x(\U891/U1118_3_/n2 ), .a(\U891/U1118_3_/n2 ), 
        .b(\U891/U1118_3_/nr ), .c(\U891/U1118_3_/nd ) );
    inv_2 \U891/U1118_3_/U3  ( .x(\a[3] ), .a(\U891/U1118_3_/n2 ) );
    nor3_1 \U891/U1117_0_/Unr  ( .x(\U891/U1117_0_/nr ), .a(i[0]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_0_/Und  ( .x(\U891/U1117_0_/nd ), .a(i[0]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_0_/U1  ( .x(\U891/U1117_0_/n2 ), .a(\U891/U1117_0_/n2 ), 
        .b(\U891/U1117_0_/nr ), .c(\U891/U1117_0_/nd ) );
    inv_2 \U891/U1117_0_/U3  ( .x(\b[0] ), .a(\U891/U1117_0_/n2 ) );
    nor3_1 \U891/U1117_1_/Unr  ( .x(\U891/U1117_1_/nr ), .a(i[1]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_1_/Und  ( .x(\U891/U1117_1_/nd ), .a(i[1]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_1_/U1  ( .x(\U891/U1117_1_/n2 ), .a(\U891/U1117_1_/n2 ), 
        .b(\U891/U1117_1_/nr ), .c(\U891/U1117_1_/nd ) );
    inv_2 \U891/U1117_1_/U3  ( .x(\b[1] ), .a(\U891/U1117_1_/n2 ) );
    nor3_1 \U891/U1117_2_/Unr  ( .x(\U891/U1117_2_/nr ), .a(i[2]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_2_/Und  ( .x(\U891/U1117_2_/nd ), .a(i[2]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_2_/U1  ( .x(\U891/U1117_2_/n2 ), .a(\U891/U1117_2_/n2 ), 
        .b(\U891/U1117_2_/nr ), .c(\U891/U1117_2_/nd ) );
    inv_2 \U891/U1117_2_/U3  ( .x(\b[2] ), .a(\U891/U1117_2_/n2 ) );
    nor3_1 \U891/U1117_3_/Unr  ( .x(\U891/U1117_3_/nr ), .a(i[3]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_3_/Und  ( .x(\U891/U1117_3_/nd ), .a(i[3]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_3_/U1  ( .x(\U891/U1117_3_/n2 ), .a(\U891/U1117_3_/n2 ), 
        .b(\U891/U1117_3_/nr ), .c(\U891/U1117_3_/nd ) );
    inv_2 \U891/U1117_3_/U3  ( .x(\b[3] ), .a(\U891/U1117_3_/n2 ) );
    inv_1 \U886/U1126/U3  ( .x(\U886/reset ), .a(nbReset) );
    nor3_1 \U886/U1128/U27  ( .x(\U886/U1128/nb ), .a(\U886/reset ), .b(\f[3] 
        ), .c(\f[2] ) );
    nor2_1 \U886/U1128/U26  ( .x(\U886/U1128/na ), .a(\f[1] ), .b(\f[0] ) );
    nand2_2 \U886/U1128/U29  ( .x(\U886/ackb ), .a(\U886/U1128/nb ), .b(
        \U886/U1128/na ) );
    nor2_1 \U886/U1108/U5  ( .x(\U886/nack ), .a(\U886/acka ), .b(\U886/ackb )
         );
    nor2_2 \U886/U914/U6  ( .x(nba), .a(\U886/acka ), .b(\U886/ackb ) );
    and4_1 \U886/U1127/U25  ( .x(\U886/U1127/n5 ), .a(\U886/U1127/n1 ), .b(
        \U886/U1127/n2 ), .c(\U886/U1127/n3 ), .d(\U886/U1127/n4 ) );
    inv_1 \U886/U1127/U1  ( .x(\U886/U1127/n1 ), .a(\e[3] ) );
    inv_1 \U886/U1127/U2  ( .x(\U886/U1127/n2 ), .a(\e[2] ) );
    inv_1 \U886/U1127/U3  ( .x(\U886/U1127/n3 ), .a(\e[1] ) );
    inv_1 \U886/U1127/U4  ( .x(\U886/U1127/n4 ), .a(\e[0] ) );
    inv_2 \U886/U1127/U5  ( .x(\U886/acka ), .a(\U886/U1127/n5 ) );
    ao222_2 \U886/U1121/U19/U1/U1  ( .x(fsela), .a(\U886/nack ), .b(fsel), .c(
        \U886/nack ), .d(fsela), .e(fsel), .f(fsela) );
    ao222_2 \U886/U1120/U19/U1/U1  ( .x(esela), .a(esel), .b(\U886/nack ), .c(
        esel), .d(esela), .e(\U886/nack ), .f(esela) );
    nor3_1 \U886/U1118_0_/Unr  ( .x(\U886/U1118_0_/nr ), .a(\b[0] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_0_/Und  ( .x(\U886/U1118_0_/nd ), .a(\b[0] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_0_/U1  ( .x(\U886/U1118_0_/n2 ), .a(\U886/U1118_0_/n2 ), 
        .b(\U886/U1118_0_/nr ), .c(\U886/U1118_0_/nd ) );
    inv_2 \U886/U1118_0_/U3  ( .x(\e[0] ), .a(\U886/U1118_0_/n2 ) );
    nor3_1 \U886/U1118_1_/Unr  ( .x(\U886/U1118_1_/nr ), .a(\b[1] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_1_/Und  ( .x(\U886/U1118_1_/nd ), .a(\b[1] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_1_/U1  ( .x(\U886/U1118_1_/n2 ), .a(\U886/U1118_1_/n2 ), 
        .b(\U886/U1118_1_/nr ), .c(\U886/U1118_1_/nd ) );
    inv_2 \U886/U1118_1_/U3  ( .x(\e[1] ), .a(\U886/U1118_1_/n2 ) );
    nor3_1 \U886/U1118_2_/Unr  ( .x(\U886/U1118_2_/nr ), .a(\b[2] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_2_/Und  ( .x(\U886/U1118_2_/nd ), .a(\b[2] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_2_/U1  ( .x(\U886/U1118_2_/n2 ), .a(\U886/U1118_2_/n2 ), 
        .b(\U886/U1118_2_/nr ), .c(\U886/U1118_2_/nd ) );
    inv_2 \U886/U1118_2_/U3  ( .x(\e[2] ), .a(\U886/U1118_2_/n2 ) );
    nor3_1 \U886/U1118_3_/Unr  ( .x(\U886/U1118_3_/nr ), .a(\b[3] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_3_/Und  ( .x(\U886/U1118_3_/nd ), .a(\b[3] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_3_/U1  ( .x(\U886/U1118_3_/n2 ), .a(\U886/U1118_3_/n2 ), 
        .b(\U886/U1118_3_/nr ), .c(\U886/U1118_3_/nd ) );
    inv_2 \U886/U1118_3_/U3  ( .x(\e[3] ), .a(\U886/U1118_3_/n2 ) );
    nor3_1 \U886/U1117_0_/Unr  ( .x(\U886/U1117_0_/nr ), .a(\b[0] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_0_/Und  ( .x(\U886/U1117_0_/nd ), .a(\b[0] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_0_/U1  ( .x(\U886/U1117_0_/n2 ), .a(\U886/U1117_0_/n2 ), 
        .b(\U886/U1117_0_/nr ), .c(\U886/U1117_0_/nd ) );
    inv_2 \U886/U1117_0_/U3  ( .x(\f[0] ), .a(\U886/U1117_0_/n2 ) );
    nor3_1 \U886/U1117_1_/Unr  ( .x(\U886/U1117_1_/nr ), .a(\b[1] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_1_/Und  ( .x(\U886/U1117_1_/nd ), .a(\b[1] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_1_/U1  ( .x(\U886/U1117_1_/n2 ), .a(\U886/U1117_1_/n2 ), 
        .b(\U886/U1117_1_/nr ), .c(\U886/U1117_1_/nd ) );
    inv_2 \U886/U1117_1_/U3  ( .x(\f[1] ), .a(\U886/U1117_1_/n2 ) );
    nor3_1 \U886/U1117_2_/Unr  ( .x(\U886/U1117_2_/nr ), .a(\b[2] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_2_/Und  ( .x(\U886/U1117_2_/nd ), .a(\b[2] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_2_/U1  ( .x(\U886/U1117_2_/n2 ), .a(\U886/U1117_2_/n2 ), 
        .b(\U886/U1117_2_/nr ), .c(\U886/U1117_2_/nd ) );
    inv_2 \U886/U1117_2_/U3  ( .x(\f[2] ), .a(\U886/U1117_2_/n2 ) );
    nor3_1 \U886/U1117_3_/Unr  ( .x(\U886/U1117_3_/nr ), .a(\b[3] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_3_/Und  ( .x(\U886/U1117_3_/nd ), .a(\b[3] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_3_/U1  ( .x(\U886/U1117_3_/n2 ), .a(\U886/U1117_3_/n2 ), 
        .b(\U886/U1117_3_/nr ), .c(\U886/U1117_3_/nd ) );
    inv_2 \U886/U1117_3_/U3  ( .x(\f[3] ), .a(\U886/U1117_3_/n2 ) );
    inv_1 \U884/U1126/U3  ( .x(\U884/reset ), .a(nbReset) );
    nor3_1 \U884/U1128/U27  ( .x(\U884/U1128/nb ), .a(\U884/reset ), .b(\d[3] 
        ), .c(\d[2] ) );
    nor2_1 \U884/U1128/U26  ( .x(\U884/U1128/na ), .a(\d[1] ), .b(\d[0] ) );
    nand2_2 \U884/U1128/U29  ( .x(\U884/ackb ), .a(\U884/U1128/nb ), .b(
        \U884/U1128/na ) );
    nor2_1 \U884/U1108/U5  ( .x(\U884/nack ), .a(\U884/acka ), .b(\U884/ackb )
         );
    nor2_2 \U884/U914/U6  ( .x(naa), .a(\U884/acka ), .b(\U884/ackb ) );
    and4_1 \U884/U1127/U25  ( .x(\U884/U1127/n5 ), .a(\U884/U1127/n1 ), .b(
        \U884/U1127/n2 ), .c(\U884/U1127/n3 ), .d(\U884/U1127/n4 ) );
    inv_1 \U884/U1127/U1  ( .x(\U884/U1127/n1 ), .a(\c[3] ) );
    inv_1 \U884/U1127/U2  ( .x(\U884/U1127/n2 ), .a(\c[2] ) );
    inv_1 \U884/U1127/U3  ( .x(\U884/U1127/n3 ), .a(\c[1] ) );
    inv_1 \U884/U1127/U4  ( .x(\U884/U1127/n4 ), .a(\c[0] ) );
    inv_2 \U884/U1127/U5  ( .x(\U884/acka ), .a(\U884/U1127/n5 ) );
    ao222_2 \U884/U1121/U19/U1/U1  ( .x(dsela), .a(\U884/nack ), .b(dsel), .c(
        \U884/nack ), .d(dsela), .e(dsel), .f(dsela) );
    ao222_2 \U884/U1120/U19/U1/U1  ( .x(csela), .a(csel), .b(\U884/nack ), .c(
        csel), .d(csela), .e(\U884/nack ), .f(csela) );
    nor3_1 \U884/U1118_0_/Unr  ( .x(\U884/U1118_0_/nr ), .a(\a[0] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_0_/Und  ( .x(\U884/U1118_0_/nd ), .a(\a[0] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_0_/U1  ( .x(\U884/U1118_0_/n2 ), .a(\U884/U1118_0_/n2 ), 
        .b(\U884/U1118_0_/nr ), .c(\U884/U1118_0_/nd ) );
    inv_2 \U884/U1118_0_/U3  ( .x(\c[0] ), .a(\U884/U1118_0_/n2 ) );
    nor3_1 \U884/U1118_1_/Unr  ( .x(\U884/U1118_1_/nr ), .a(\a[1] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_1_/Und  ( .x(\U884/U1118_1_/nd ), .a(\a[1] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_1_/U1  ( .x(\U884/U1118_1_/n2 ), .a(\U884/U1118_1_/n2 ), 
        .b(\U884/U1118_1_/nr ), .c(\U884/U1118_1_/nd ) );
    inv_2 \U884/U1118_1_/U3  ( .x(\c[1] ), .a(\U884/U1118_1_/n2 ) );
    nor3_1 \U884/U1118_2_/Unr  ( .x(\U884/U1118_2_/nr ), .a(\a[2] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_2_/Und  ( .x(\U884/U1118_2_/nd ), .a(\a[2] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_2_/U1  ( .x(\U884/U1118_2_/n2 ), .a(\U884/U1118_2_/n2 ), 
        .b(\U884/U1118_2_/nr ), .c(\U884/U1118_2_/nd ) );
    inv_2 \U884/U1118_2_/U3  ( .x(\c[2] ), .a(\U884/U1118_2_/n2 ) );
    nor3_1 \U884/U1118_3_/Unr  ( .x(\U884/U1118_3_/nr ), .a(\a[3] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_3_/Und  ( .x(\U884/U1118_3_/nd ), .a(\a[3] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_3_/U1  ( .x(\U884/U1118_3_/n2 ), .a(\U884/U1118_3_/n2 ), 
        .b(\U884/U1118_3_/nr ), .c(\U884/U1118_3_/nd ) );
    inv_2 \U884/U1118_3_/U3  ( .x(\c[3] ), .a(\U884/U1118_3_/n2 ) );
    nor3_1 \U884/U1117_0_/Unr  ( .x(\U884/U1117_0_/nr ), .a(\a[0] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_0_/Und  ( .x(\U884/U1117_0_/nd ), .a(\a[0] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_0_/U1  ( .x(\U884/U1117_0_/n2 ), .a(\U884/U1117_0_/n2 ), 
        .b(\U884/U1117_0_/nr ), .c(\U884/U1117_0_/nd ) );
    inv_2 \U884/U1117_0_/U3  ( .x(\d[0] ), .a(\U884/U1117_0_/n2 ) );
    nor3_1 \U884/U1117_1_/Unr  ( .x(\U884/U1117_1_/nr ), .a(\a[1] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_1_/Und  ( .x(\U884/U1117_1_/nd ), .a(\a[1] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_1_/U1  ( .x(\U884/U1117_1_/n2 ), .a(\U884/U1117_1_/n2 ), 
        .b(\U884/U1117_1_/nr ), .c(\U884/U1117_1_/nd ) );
    inv_2 \U884/U1117_1_/U3  ( .x(\d[1] ), .a(\U884/U1117_1_/n2 ) );
    nor3_1 \U884/U1117_2_/Unr  ( .x(\U884/U1117_2_/nr ), .a(\a[2] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_2_/Und  ( .x(\U884/U1117_2_/nd ), .a(\a[2] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_2_/U1  ( .x(\U884/U1117_2_/n2 ), .a(\U884/U1117_2_/n2 ), 
        .b(\U884/U1117_2_/nr ), .c(\U884/U1117_2_/nd ) );
    inv_2 \U884/U1117_2_/U3  ( .x(\d[2] ), .a(\U884/U1117_2_/n2 ) );
    nor3_1 \U884/U1117_3_/Unr  ( .x(\U884/U1117_3_/nr ), .a(\a[3] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_3_/Und  ( .x(\U884/U1117_3_/nd ), .a(\a[3] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_3_/U1  ( .x(\U884/U1117_3_/n2 ), .a(\U884/U1117_3_/n2 ), 
        .b(\U884/U1117_3_/nr ), .c(\U884/U1117_3_/nd ) );
    inv_2 \U884/U1117_3_/U3  ( .x(\d[3] ), .a(\U884/U1117_3_/n2 ) );
    nand2_1 \U888/U1128/U5  ( .x(\U888/s ), .a(\U888/r ), .b(\U888/nback ) );
    nand2_1 \U888/U1103/U5  ( .x(\U888/r ), .a(\U888/naack ), .b(\U888/s ) );
    inv_1 \U888/U1111/U3  ( .x(\U888/reset ), .a(nbReset) );
    inv_1 \U888/U1112/U3  ( .x(\U888/naack ), .a(esela) );
    nor2_1 \U888/U1127/U5  ( .x(\U888/nback ), .a(fsela), .b(\U888/reset ) );
    and2_2 \U888/U1129/U8  ( .x(esel), .a(\U888/nback ), .b(\U888/s ) );
    and2_2 \U888/U1124/U8  ( .x(fsel), .a(\U888/r ), .b(\U888/naack ) );
    nand2_1 \U887/U1128/U5  ( .x(\U887/s ), .a(\U887/r ), .b(\U887/nback ) );
    nand2_1 \U887/U1103/U5  ( .x(\U887/r ), .a(\U887/naack ), .b(\U887/s ) );
    inv_1 \U887/U1111/U3  ( .x(\U887/reset ), .a(nbReset) );
    inv_1 \U887/U1112/U3  ( .x(\U887/naack ), .a(csela) );
    nor2_1 \U887/U1127/U5  ( .x(\U887/nback ), .a(dsela), .b(\U887/reset ) );
    and2_2 \U887/U1129/U8  ( .x(csel), .a(\U887/nback ), .b(\U887/s ) );
    and2_2 \U887/U1124/U8  ( .x(dsel), .a(\U887/r ), .b(\U887/naack ) );
    nand2_1 \U885/U1128/U5  ( .x(\U885/s ), .a(\U885/r ), .b(\U885/nback ) );
    nand2_1 \U885/U1103/U5  ( .x(\U885/r ), .a(\U885/naack ), .b(\U885/s ) );
    inv_1 \U885/U1111/U3  ( .x(\U885/reset ), .a(nbReset) );
    inv_1 \U885/U1112/U3  ( .x(\U885/naack ), .a(asela) );
    nor2_1 \U885/U1127/U5  ( .x(\U885/nback ), .a(bsela), .b(\U885/reset ) );
    and2_2 \U885/U1129/U8  ( .x(asel), .a(\U885/nback ), .b(\U885/s ) );
    and2_2 \U885/U1124/U8  ( .x(bsel), .a(\U885/r ), .b(\U885/naack ) );
    nor3_1 \U877/U594/U7  ( .x(\U877/x ), .a(ol[7]), .b(\U877/reset ), .c(oh
        [7]) );
    nor3_1 \U877/U593/U7  ( .x(\U877/y ), .a(ol[6]), .b(\U877/reset ), .c(oh
        [6]) );
    inv_1 \U877/U604/U3  ( .x(\U877/reset ), .a(nbReset) );
    oa31_1 \U877/U590/U25/U1/Uclr  ( .x(\U877/U590/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[1] ), .d(oh[6]) );
    oaoi211_1 \U877/U590/U25/U1/Uaoi  ( .x(\U877/U590/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[1] ), .c(n1), .d(\U877/U590/U25/U1/clr ) );
    inv_2 \U877/U590/U25/U1/Ui  ( .x(oh[6]), .a(\U877/U590/U25/U1/ob ) );
    oa31_1 \U877/U589/U25/U1/Uclr  ( .x(\U877/U589/U25/U1/clr ), .a(net135), 
        .b(\cl[1] ), .c(\cl[0] ), .d(ol[7]) );
    oaoi211_1 \U877/U589/U25/U1/Uaoi  ( .x(\U877/U589/U25/U1/ob ), .a(\cl[1] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U589/U25/U1/clr ) );
    inv_2 \U877/U589/U25/U1/Ui  ( .x(ol[7]), .a(\U877/U589/U25/U1/ob ) );
    oa31_1 \U877/U588/U25/U1/Uclr  ( .x(\U877/U588/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[2] ), .d(oh[7]) );
    oaoi211_1 \U877/U588/U25/U1/Uaoi  ( .x(\U877/U588/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[2] ), .c(n1), .d(\U877/U588/U25/U1/clr ) );
    inv_2 \U877/U588/U25/U1/Ui  ( .x(oh[7]), .a(\U877/U588/U25/U1/ob ) );
    oa31_1 \U877/U591/U25/U1/Uclr  ( .x(\U877/U591/U25/U1/clr ), .a(net135), 
        .b(\cl[2] ), .c(\cl[0] ), .d(ol[6]) );
    oaoi211_1 \U877/U591/U25/U1/Uaoi  ( .x(\U877/U591/U25/U1/ob ), .a(\cl[2] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U591/U25/U1/clr ) );
    inv_2 \U877/U591/U25/U1/Ui  ( .x(ol[6]), .a(\U877/U591/U25/U1/ob ) );
    ao222_2 \U877/U592/U19/U1/U1  ( .x(ncla), .a(\U877/x ), .b(\U877/y ), .c(
        \U877/x ), .d(ncla), .e(\U877/y ), .f(ncla) );
    nor3_1 \U876/U594/U7  ( .x(\U876/x ), .a(ol[3]), .b(\U876/reset ), .c(oh
        [3]) );
    nor3_1 \U876/U593/U7  ( .x(\U876/y ), .a(ol[2]), .b(\U876/reset ), .c(oh
        [2]) );
    inv_1 \U876/U604/U3  ( .x(\U876/reset ), .a(nbReset) );
    oa31_1 \U876/U590/U25/U1/Uclr  ( .x(\U876/U590/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[1] ), .d(oh[2]) );
    oaoi211_1 \U876/U590/U25/U1/Uaoi  ( .x(\U876/U590/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[1] ), .c(n1), .d(\U876/U590/U25/U1/clr ) );
    inv_2 \U876/U590/U25/U1/Ui  ( .x(oh[2]), .a(\U876/U590/U25/U1/ob ) );
    oa31_1 \U876/U589/U25/U1/Uclr  ( .x(\U876/U589/U25/U1/clr ), .a(net135), 
        .b(\d[1] ), .c(\d[0] ), .d(ol[3]) );
    oaoi211_1 \U876/U589/U25/U1/Uaoi  ( .x(\U876/U589/U25/U1/ob ), .a(\d[1] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U589/U25/U1/clr ) );
    inv_2 \U876/U589/U25/U1/Ui  ( .x(ol[3]), .a(\U876/U589/U25/U1/ob ) );
    oa31_1 \U876/U588/U25/U1/Uclr  ( .x(\U876/U588/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[2] ), .d(oh[3]) );
    oaoi211_1 \U876/U588/U25/U1/Uaoi  ( .x(\U876/U588/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[2] ), .c(n1), .d(\U876/U588/U25/U1/clr ) );
    inv_2 \U876/U588/U25/U1/Ui  ( .x(oh[3]), .a(\U876/U588/U25/U1/ob ) );
    oa31_1 \U876/U591/U25/U1/Uclr  ( .x(\U876/U591/U25/U1/clr ), .a(net135), 
        .b(\d[2] ), .c(\d[0] ), .d(ol[2]) );
    oaoi211_1 \U876/U591/U25/U1/Uaoi  ( .x(\U876/U591/U25/U1/ob ), .a(\d[2] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U591/U25/U1/clr ) );
    inv_2 \U876/U591/U25/U1/Ui  ( .x(ol[2]), .a(\U876/U591/U25/U1/ob ) );
    ao222_2 \U876/U592/U19/U1/U1  ( .x(nda), .a(\U876/x ), .b(\U876/y ), .c(
        \U876/x ), .d(nda), .e(\U876/y ), .f(nda) );
    nor3_1 \U2/U594/U7  ( .x(\U2/x ), .a(ol[1]), .b(\U2/reset ), .c(oh[1]) );
    nor3_1 \U2/U593/U7  ( .x(\U2/y ), .a(ol[0]), .b(\U2/reset ), .c(oh[0]) );
    inv_1 \U2/U604/U3  ( .x(\U2/reset ), .a(nbReset) );
    oa31_1 \U2/U590/U25/U1/Uclr  ( .x(\U2/U590/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[1] ), .d(oh[0]) );
    oaoi211_1 \U2/U590/U25/U1/Uaoi  ( .x(\U2/U590/U25/U1/ob ), .a(\f[3] ), .b(
        \f[1] ), .c(n1), .d(\U2/U590/U25/U1/clr ) );
    inv_2 \U2/U590/U25/U1/Ui  ( .x(oh[0]), .a(\U2/U590/U25/U1/ob ) );
    oa31_1 \U2/U589/U25/U1/Uclr  ( .x(\U2/U589/U25/U1/clr ), .a(net135), .b(
        \f[1] ), .c(\f[0] ), .d(ol[1]) );
    oaoi211_1 \U2/U589/U25/U1/Uaoi  ( .x(\U2/U589/U25/U1/ob ), .a(\f[1] ), .b(
        \f[0] ), .c(n1), .d(\U2/U589/U25/U1/clr ) );
    inv_2 \U2/U589/U25/U1/Ui  ( .x(ol[1]), .a(\U2/U589/U25/U1/ob ) );
    oa31_1 \U2/U588/U25/U1/Uclr  ( .x(\U2/U588/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[2] ), .d(oh[1]) );
    oaoi211_1 \U2/U588/U25/U1/Uaoi  ( .x(\U2/U588/U25/U1/ob ), .a(\f[3] ), .b(
        \f[2] ), .c(n1), .d(\U2/U588/U25/U1/clr ) );
    inv_2 \U2/U588/U25/U1/Ui  ( .x(oh[1]), .a(\U2/U588/U25/U1/ob ) );
    oa31_1 \U2/U591/U25/U1/Uclr  ( .x(\U2/U591/U25/U1/clr ), .a(net135), .b(
        \f[2] ), .c(\f[0] ), .d(ol[0]) );
    oaoi211_1 \U2/U591/U25/U1/Uaoi  ( .x(\U2/U591/U25/U1/ob ), .a(\f[2] ), .b(
        \f[0] ), .c(n1), .d(\U2/U591/U25/U1/clr ) );
    inv_2 \U2/U591/U25/U1/Ui  ( .x(ol[0]), .a(\U2/U591/U25/U1/ob ) );
    ao222_2 \U2/U592/U19/U1/U1  ( .x(nfa), .a(\U2/x ), .b(\U2/y ), .c(\U2/x ), 
        .d(nfa), .e(\U2/y ), .f(nfa) );
    nor3_1 \U1/U594/U7  ( .x(\U1/x ), .a(ol[5]), .b(\U1/reset ), .c(oh[5]) );
    nor3_1 \U1/U593/U7  ( .x(\U1/y ), .a(ol[4]), .b(\U1/reset ), .c(oh[4]) );
    inv_1 \U1/U604/U3  ( .x(\U1/reset ), .a(nbReset) );
    oa31_1 \U1/U590/U25/U1/Uclr  ( .x(\U1/U590/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[1] ), .d(oh[4]) );
    oaoi211_1 \U1/U590/U25/U1/Uaoi  ( .x(\U1/U590/U25/U1/ob ), .a(\e[3] ), .b(
        \e[1] ), .c(n1), .d(\U1/U590/U25/U1/clr ) );
    inv_2 \U1/U590/U25/U1/Ui  ( .x(oh[4]), .a(\U1/U590/U25/U1/ob ) );
    oa31_1 \U1/U589/U25/U1/Uclr  ( .x(\U1/U589/U25/U1/clr ), .a(net135), .b(
        \e[1] ), .c(\e[0] ), .d(ol[5]) );
    oaoi211_1 \U1/U589/U25/U1/Uaoi  ( .x(\U1/U589/U25/U1/ob ), .a(\e[1] ), .b(
        \e[0] ), .c(n1), .d(\U1/U589/U25/U1/clr ) );
    inv_2 \U1/U589/U25/U1/Ui  ( .x(ol[5]), .a(\U1/U589/U25/U1/ob ) );
    oa31_1 \U1/U588/U25/U1/Uclr  ( .x(\U1/U588/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[2] ), .d(oh[5]) );
    oaoi211_1 \U1/U588/U25/U1/Uaoi  ( .x(\U1/U588/U25/U1/ob ), .a(\e[3] ), .b(
        \e[2] ), .c(n1), .d(\U1/U588/U25/U1/clr ) );
    inv_2 \U1/U588/U25/U1/Ui  ( .x(oh[5]), .a(\U1/U588/U25/U1/ob ) );
    oa31_1 \U1/U591/U25/U1/Uclr  ( .x(\U1/U591/U25/U1/clr ), .a(net135), .b(
        \e[2] ), .c(\e[0] ), .d(ol[4]) );
    oaoi211_1 \U1/U591/U25/U1/Uaoi  ( .x(\U1/U591/U25/U1/ob ), .a(\e[2] ), .b(
        \e[0] ), .c(n1), .d(\U1/U591/U25/U1/clr ) );
    inv_2 \U1/U591/U25/U1/Ui  ( .x(ol[4]), .a(\U1/U591/U25/U1/ob ) );
    ao222_2 \U1/U592/U19/U1/U1  ( .x(nea), .a(\U1/x ), .b(\U1/y ), .c(\U1/x ), 
        .d(nea), .e(\U1/y ), .f(nea) );
    and3_4 \U881/U20/U9  ( .x(nca), .a(\U881/nack[1] ), .b(\U881/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U881/U18/U5  ( .x(\U881/nack[0] ), .a(\cl[3] ), .b(\cl[0] ) );
    nor2_1 \U881/U19/U5  ( .x(\U881/nack[1] ), .a(\cl[1] ), .b(\cl[2] ) );
    ao222_2 \U881/U15_0_/U19/U1/U1  ( .x(\cl[0] ), .a(\c[0] ), .b(ncla), .c(
        \c[0] ), .d(\cl[0] ), .e(ncla), .f(\cl[0] ) );
    ao222_2 \U881/U15_1_/U19/U1/U1  ( .x(\cl[1] ), .a(\c[1] ), .b(ncla), .c(
        \c[1] ), .d(\cl[1] ), .e(ncla), .f(\cl[1] ) );
    ao222_2 \U881/U15_2_/U19/U1/U1  ( .x(\cl[2] ), .a(\c[2] ), .b(ncla), .c(
        \c[2] ), .d(\cl[2] ), .e(ncla), .f(\cl[2] ) );
    ao222_2 \U881/U15_3_/U19/U1/U1  ( .x(\cl[3] ), .a(\c[3] ), .b(ncla), .c(
        \c[3] ), .d(\cl[3] ), .e(ncla), .f(\cl[3] ) );
    and2_5 U1 ( .x(n1), .a(nbReset), .b(noa) );
    and2_3 U2 ( .x(net135), .a(nbReset), .b(noa) );
endmodule


module chain_dr2fr_byte_1 ( eop_ack, ia, o, eop, ih, il, nReset, noa );
output [4:0] o;
input  [7:0] ih;
input  [7:0] il;
input  eop, nReset, noa;
output eop_ack, ia;
    wire eop_pass, nhighack, nlowack, \twobitack[2] , \twobitack[3] , 
        \twobitack[0] , \twobitack[1] , xsel, ysel, nxa, nyla, nbReset, nya, 
        \y[3] , \y[2] , \y[1] , \y[0] , \yl[3] , \yl[2] , \yl[1] , \yl[0] , 
        \cdh[0] , \cdh[1] , \cdl[0] , \cdl[1] , net193, \cdh[2] , \cdh[3] , 
        \cdl[2] , \cdl[3] , net195, bsel, dsel, nba, bg, nda, dg, asel, csel, 
        naa, ag, nca, cg, \d[3] , \d[2] , \d[1] , \d[0] , \b[3] , \b[2] , 
        \b[1] , \b[0] , \x[3] , \x[2] , \x[1] , \x[0] , \c[3] , \c[2] , \c[1] , 
        \c[0] , \a[3] , \a[2] , \a[1] , \a[0] , net194, net199, \U1018/Z , 
        \U1270/net190 , \U1270/net191 , \U1270/net192 , \U1270/net189 , 
        \U1270/U1141/Z , \U1268/net190 , \U1268/net191 , \U1268/net192 , 
        \U1268/net189 , \U1268/U1141/Z , \U1224/nack[0] , \U1224/nack[1] , 
        \U1224/net4 , \U1224/U1125/U28/U1/clr , \U1224/U1125/U28/U1/set , 
        \U1224/U1122/U28/U1/clr , \U1224/U1122/U28/U1/set , 
        \U1224/U916_0_/U25/U1/clr , \U1224/U916_0_/U25/U1/ob , 
        \U1224/U916_1_/U25/U1/clr , \U1224/U916_1_/U25/U1/ob , 
        \U1224/U916_2_/U25/U1/clr , \U1224/U916_2_/U25/U1/ob , 
        \U1224/U916_3_/U25/U1/clr , \U1224/U916_3_/U25/U1/ob , \U1209/nack[0] , 
        \U1209/nack[1] , \U1209/net4 , \U1209/U1125/U28/U1/clr , 
        \U1209/U1125/U28/U1/set , \U1209/U1122/U28/U1/clr , 
        \U1209/U1122/U28/U1/set , \U1209/U916_0_/U25/U1/clr , 
        \U1209/U916_0_/U25/U1/ob , \U1209/U916_1_/U25/U1/clr , 
        \U1209/U916_1_/U25/U1/ob , \U1209/U916_2_/U25/U1/clr , 
        \U1209/U916_2_/U25/U1/ob , \U1209/U916_3_/U25/U1/clr , 
        \U1209/U916_3_/U25/U1/ob , \U1213/nack[0] , \U1213/nack[1] , 
        \U1213/net4 , \U1213/U1125/U28/U1/clr , \U1213/U1125/U28/U1/set , 
        \U1213/U1122/U28/U1/clr , \U1213/U1122/U28/U1/set , 
        \U1213/U916_0_/U25/U1/clr , \U1213/U916_0_/U25/U1/ob , 
        \U1213/U916_1_/U25/U1/clr , \U1213/U916_1_/U25/U1/ob , 
        \U1213/U916_2_/U25/U1/clr , \U1213/U916_2_/U25/U1/ob , 
        \U1213/U916_3_/U25/U1/clr , \U1213/U916_3_/U25/U1/ob , \U1296/ng , 
        \U1296/U1384/Z , \U1296/U1386/U25/U1/clr , \U1296/U1386/U25/U1/ob , 
        \U1298/ng , \U1298/U1384/Z , \U1298/U1386/U25/U1/clr , 
        \U1298/U1386/U25/U1/ob , \U1306/ng , \U1306/U1384/Z , 
        \U1306/U1386/U25/U1/clr , \U1306/U1386/U25/U1/ob , \U1295/ng , 
        \U1295/U1384/Z , \U1295/U1386/U25/U1/clr , \U1295/U1386/U25/U1/ob , 
        \U1297/s , \U1297/nback , \U1297/r , \U1297/naack , \U1297/reset , 
        \U1297/U1128/U28/U1/clr , \U1297/U1128/U28/U1/set , 
        \U1297/U1127/U28/U1/clr , \U1297/U1127/U28/U1/set , \U1300/s , 
        \U1300/nback , \U1300/r , \U1300/naack , \U1300/reset , 
        \U1300/U1128/U28/U1/clr , \U1300/U1128/U28/U1/set , 
        \U1300/U1127/U28/U1/clr , \U1300/U1127/U28/U1/set , \U1289/bnreset , 
        \U1289/U1150/U28/U1/clr , \U1289/U1150/U28/U1/set , 
        \U1289/U1152/U28/U1/clr , \U1289/U1152/U28/U1/set , 
        \U1289/U1149/U28/U1/clr , \U1289/U1149/U28/U1/set , 
        \U1289/U1151/U28/U1/clr , \U1289/U1151/U28/U1/set , 
        \U1289/U1148/net190 , \U1289/U1148/net191 , \U1289/U1148/net192 , 
        \U1289/U1148/net189 , \U1289/U1148/U1141/Z , \U1271/bnreset , 
        \U1271/U1150/U28/U1/clr , \U1271/U1150/U28/U1/set , 
        \U1271/U1152/U28/U1/clr , \U1271/U1152/U28/U1/set , 
        \U1271/U1149/U28/U1/clr , \U1271/U1149/U28/U1/set , 
        \U1271/U1151/U28/U1/clr , \U1271/U1151/U28/U1/set , 
        \U1271/U1148/net190 , \U1271/U1148/net191 , \U1271/U1148/net192 , 
        \U1271/U1148/net189 , \U1271/U1148/U1141/Z , \U1225/naack , \U1225/r , 
        \U1225/s , \U1225/nback , \U1225/reset , \U1308/nack[1] , 
        \U1308/nack[0] ;
    assign o[4] = eop_ack;
    buf_2 U1231 ( .x(nbReset), .a(nReset) );
    and3_1 \U1194/U9  ( .x(eop_pass), .a(nxa), .b(naa), .c(eop) );
    ao222_1 \U1301/U18/U1/U1  ( .x(nlowack), .a(\twobitack[0] ), .b(
        \twobitack[1] ), .c(\twobitack[0] ), .d(nlowack), .e(\twobitack[1] ), 
        .f(nlowack) );
    ao222_1 \U1302/U18/U1/U1  ( .x(nhighack), .a(\twobitack[2] ), .b(
        \twobitack[3] ), .c(\twobitack[2] ), .d(nhighack), .e(\twobitack[3] ), 
        .f(nhighack) );
    aoi222_1 \U1018/U30/U1  ( .x(ia), .a(nhighack), .b(nlowack), .c(nhighack), 
        .d(\U1018/Z ), .e(nlowack), .f(\U1018/Z ) );
    inv_1 \U1018/U30/Uinv  ( .x(\U1018/Z ), .a(ia) );
    ao222_2 \U1038/U19/U1/U1  ( .x(eop_ack), .a(eop_pass), .b(noa), .c(
        eop_pass), .d(eop_ack), .e(noa), .f(eop_ack) );
    inv_1 \U1270/U1147/U3  ( .x(\U1270/net189 ), .a(nbReset) );
    nor2_1 \U1270/U582/U5  ( .x(\U1270/net192 ), .a(il[4]), .b(ih[4]) );
    nor2_1 \U1270/U580/U5  ( .x(\U1270/net191 ), .a(il[5]), .b(ih[5]) );
    nor2_2 \U1270/U1146/U6  ( .x(net199), .a(\U1270/net190 ), .b(
        \U1270/net189 ) );
    aoi222_1 \U1270/U1141/U30/U1  ( .x(\U1270/net190 ), .a(\U1270/net191 ), 
        .b(\U1270/net192 ), .c(\U1270/net191 ), .d(\U1270/U1141/Z ), .e(
        \U1270/net192 ), .f(\U1270/U1141/Z ) );
    inv_1 \U1270/U1141/U30/Uinv  ( .x(\U1270/U1141/Z ), .a(\U1270/net190 ) );
    inv_1 \U1268/U1147/U3  ( .x(\U1268/net189 ), .a(nbReset) );
    nor2_1 \U1268/U582/U5  ( .x(\U1268/net192 ), .a(il[6]), .b(ih[6]) );
    nor2_1 \U1268/U580/U5  ( .x(\U1268/net191 ), .a(il[7]), .b(ih[7]) );
    nor2_2 \U1268/U1146/U6  ( .x(net194), .a(\U1268/net190 ), .b(
        \U1268/net189 ) );
    aoi222_1 \U1268/U1141/U30/U1  ( .x(\U1268/net190 ), .a(\U1268/net191 ), 
        .b(\U1268/net192 ), .c(\U1268/net191 ), .d(\U1268/U1141/Z ), .e(
        \U1268/net192 ), .f(\U1268/U1141/Z ) );
    inv_1 \U1268/U1141/U30/Uinv  ( .x(\U1268/U1141/Z ), .a(\U1268/net190 ) );
    nor2_1 \U1224/U1128/U5  ( .x(\U1224/nack[0] ), .a(\x[3] ), .b(\x[2] ) );
    nor3_1 \U1224/U1127/U7  ( .x(\U1224/nack[1] ), .a(\x[1] ), .b(\U1224/net4 
        ), .c(\x[0] ) );
    inv_1 \U1224/U907/U3  ( .x(\U1224/net4 ), .a(nbReset) );
    aoai211_1 \U1224/U1125/U28/U1/U1  ( .x(\U1224/U1125/U28/U1/clr ), .a(
        \U1224/nack[1] ), .b(\U1224/nack[0] ), .c(asel), .d(naa) );
    nand3_1 \U1224/U1125/U28/U1/U2  ( .x(\U1224/U1125/U28/U1/set ), .a(asel), 
        .b(\U1224/nack[1] ), .c(\U1224/nack[0] ) );
    nand2_2 \U1224/U1125/U28/U1/U3  ( .x(naa), .a(\U1224/U1125/U28/U1/clr ), 
        .b(\U1224/U1125/U28/U1/set ) );
    aoai211_1 \U1224/U1122/U28/U1/U1  ( .x(\U1224/U1122/U28/U1/clr ), .a(
        \U1224/nack[0] ), .b(\U1224/nack[1] ), .c(csel), .d(nca) );
    nand3_1 \U1224/U1122/U28/U1/U2  ( .x(\U1224/U1122/U28/U1/set ), .a(csel), 
        .b(\U1224/nack[0] ), .c(\U1224/nack[1] ) );
    nand2_2 \U1224/U1122/U28/U1/U3  ( .x(nca), .a(\U1224/U1122/U28/U1/clr ), 
        .b(\U1224/U1122/U28/U1/set ) );
    oa31_1 \U1224/U916_0_/U25/U1/Uclr  ( .x(\U1224/U916_0_/U25/U1/clr ), .a(
        nxa), .b(\a[0] ), .c(\c[0] ), .d(\x[0] ) );
    oaoi211_1 \U1224/U916_0_/U25/U1/Uaoi  ( .x(\U1224/U916_0_/U25/U1/ob ), .a(
        \a[0] ), .b(\c[0] ), .c(nxa), .d(\U1224/U916_0_/U25/U1/clr ) );
    inv_2 \U1224/U916_0_/U25/U1/Ui  ( .x(\x[0] ), .a(\U1224/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_1_/U25/U1/Uclr  ( .x(\U1224/U916_1_/U25/U1/clr ), .a(
        nxa), .b(\a[1] ), .c(\c[1] ), .d(\x[1] ) );
    oaoi211_1 \U1224/U916_1_/U25/U1/Uaoi  ( .x(\U1224/U916_1_/U25/U1/ob ), .a(
        \a[1] ), .b(\c[1] ), .c(nxa), .d(\U1224/U916_1_/U25/U1/clr ) );
    inv_2 \U1224/U916_1_/U25/U1/Ui  ( .x(\x[1] ), .a(\U1224/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_2_/U25/U1/Uclr  ( .x(\U1224/U916_2_/U25/U1/clr ), .a(
        nxa), .b(\a[2] ), .c(\c[2] ), .d(\x[2] ) );
    oaoi211_1 \U1224/U916_2_/U25/U1/Uaoi  ( .x(\U1224/U916_2_/U25/U1/ob ), .a(
        \a[2] ), .b(\c[2] ), .c(nxa), .d(\U1224/U916_2_/U25/U1/clr ) );
    inv_2 \U1224/U916_2_/U25/U1/Ui  ( .x(\x[2] ), .a(\U1224/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_3_/U25/U1/Uclr  ( .x(\U1224/U916_3_/U25/U1/clr ), .a(
        nxa), .b(\a[3] ), .c(\c[3] ), .d(\x[3] ) );
    oaoi211_1 \U1224/U916_3_/U25/U1/Uaoi  ( .x(\U1224/U916_3_/U25/U1/ob ), .a(
        \a[3] ), .b(\c[3] ), .c(nxa), .d(\U1224/U916_3_/U25/U1/clr ) );
    inv_2 \U1224/U916_3_/U25/U1/Ui  ( .x(\x[3] ), .a(\U1224/U916_3_/U25/U1/ob 
        ) );
    nor2_1 \U1209/U1128/U5  ( .x(\U1209/nack[0] ), .a(o[3]), .b(o[2]) );
    nor3_1 \U1209/U1127/U7  ( .x(\U1209/nack[1] ), .a(o[1]), .b(\U1209/net4 ), 
        .c(o[0]) );
    inv_1 \U1209/U907/U3  ( .x(\U1209/net4 ), .a(nbReset) );
    aoai211_1 \U1209/U1125/U28/U1/U1  ( .x(\U1209/U1125/U28/U1/clr ), .a(
        \U1209/nack[1] ), .b(\U1209/nack[0] ), .c(xsel), .d(nxa) );
    nand3_1 \U1209/U1125/U28/U1/U2  ( .x(\U1209/U1125/U28/U1/set ), .a(xsel), 
        .b(\U1209/nack[1] ), .c(\U1209/nack[0] ) );
    nand2_2 \U1209/U1125/U28/U1/U3  ( .x(nxa), .a(\U1209/U1125/U28/U1/clr ), 
        .b(\U1209/U1125/U28/U1/set ) );
    aoai211_1 \U1209/U1122/U28/U1/U1  ( .x(\U1209/U1122/U28/U1/clr ), .a(
        \U1209/nack[0] ), .b(\U1209/nack[1] ), .c(ysel), .d(nyla) );
    nand3_1 \U1209/U1122/U28/U1/U2  ( .x(\U1209/U1122/U28/U1/set ), .a(ysel), 
        .b(\U1209/nack[0] ), .c(\U1209/nack[1] ) );
    nand2_2 \U1209/U1122/U28/U1/U3  ( .x(nyla), .a(\U1209/U1122/U28/U1/clr ), 
        .b(\U1209/U1122/U28/U1/set ) );
    oa31_1 \U1209/U916_0_/U25/U1/Uclr  ( .x(\U1209/U916_0_/U25/U1/clr ), .a(
        noa), .b(\x[0] ), .c(\yl[0] ), .d(o[0]) );
    oaoi211_1 \U1209/U916_0_/U25/U1/Uaoi  ( .x(\U1209/U916_0_/U25/U1/ob ), .a(
        \x[0] ), .b(\yl[0] ), .c(noa), .d(\U1209/U916_0_/U25/U1/clr ) );
    inv_2 \U1209/U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U1209/U916_0_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_1_/U25/U1/Uclr  ( .x(\U1209/U916_1_/U25/U1/clr ), .a(
        noa), .b(\x[1] ), .c(\yl[1] ), .d(o[1]) );
    oaoi211_1 \U1209/U916_1_/U25/U1/Uaoi  ( .x(\U1209/U916_1_/U25/U1/ob ), .a(
        \x[1] ), .b(\yl[1] ), .c(noa), .d(\U1209/U916_1_/U25/U1/clr ) );
    inv_2 \U1209/U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U1209/U916_1_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_2_/U25/U1/Uclr  ( .x(\U1209/U916_2_/U25/U1/clr ), .a(
        noa), .b(\x[2] ), .c(\yl[2] ), .d(o[2]) );
    oaoi211_1 \U1209/U916_2_/U25/U1/Uaoi  ( .x(\U1209/U916_2_/U25/U1/ob ), .a(
        \x[2] ), .b(\yl[2] ), .c(noa), .d(\U1209/U916_2_/U25/U1/clr ) );
    inv_2 \U1209/U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U1209/U916_2_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_3_/U25/U1/Uclr  ( .x(\U1209/U916_3_/U25/U1/clr ), .a(
        noa), .b(\x[3] ), .c(\yl[3] ), .d(o[3]) );
    oaoi211_1 \U1209/U916_3_/U25/U1/Uaoi  ( .x(\U1209/U916_3_/U25/U1/ob ), .a(
        \x[3] ), .b(\yl[3] ), .c(noa), .d(\U1209/U916_3_/U25/U1/clr ) );
    inv_2 \U1209/U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U1209/U916_3_/U25/U1/ob )
         );
    nor2_1 \U1213/U1128/U5  ( .x(\U1213/nack[0] ), .a(\y[3] ), .b(\y[2] ) );
    nor3_1 \U1213/U1127/U7  ( .x(\U1213/nack[1] ), .a(\y[1] ), .b(\U1213/net4 
        ), .c(\y[0] ) );
    inv_1 \U1213/U907/U3  ( .x(\U1213/net4 ), .a(nbReset) );
    aoai211_1 \U1213/U1125/U28/U1/U1  ( .x(\U1213/U1125/U28/U1/clr ), .a(
        \U1213/nack[1] ), .b(\U1213/nack[0] ), .c(bsel), .d(nba) );
    nand3_1 \U1213/U1125/U28/U1/U2  ( .x(\U1213/U1125/U28/U1/set ), .a(bsel), 
        .b(\U1213/nack[1] ), .c(\U1213/nack[0] ) );
    nand2_2 \U1213/U1125/U28/U1/U3  ( .x(nba), .a(\U1213/U1125/U28/U1/clr ), 
        .b(\U1213/U1125/U28/U1/set ) );
    aoai211_1 \U1213/U1122/U28/U1/U1  ( .x(\U1213/U1122/U28/U1/clr ), .a(
        \U1213/nack[0] ), .b(\U1213/nack[1] ), .c(dsel), .d(nda) );
    nand3_1 \U1213/U1122/U28/U1/U2  ( .x(\U1213/U1122/U28/U1/set ), .a(dsel), 
        .b(\U1213/nack[0] ), .c(\U1213/nack[1] ) );
    nand2_2 \U1213/U1122/U28/U1/U3  ( .x(nda), .a(\U1213/U1122/U28/U1/clr ), 
        .b(\U1213/U1122/U28/U1/set ) );
    oa31_1 \U1213/U916_0_/U25/U1/Uclr  ( .x(\U1213/U916_0_/U25/U1/clr ), .a(
        nya), .b(\b[0] ), .c(\d[0] ), .d(\y[0] ) );
    oaoi211_1 \U1213/U916_0_/U25/U1/Uaoi  ( .x(\U1213/U916_0_/U25/U1/ob ), .a(
        \b[0] ), .b(\d[0] ), .c(nya), .d(\U1213/U916_0_/U25/U1/clr ) );
    inv_2 \U1213/U916_0_/U25/U1/Ui  ( .x(\y[0] ), .a(\U1213/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_1_/U25/U1/Uclr  ( .x(\U1213/U916_1_/U25/U1/clr ), .a(
        nya), .b(\b[1] ), .c(\d[1] ), .d(\y[1] ) );
    oaoi211_1 \U1213/U916_1_/U25/U1/Uaoi  ( .x(\U1213/U916_1_/U25/U1/ob ), .a(
        \b[1] ), .b(\d[1] ), .c(nya), .d(\U1213/U916_1_/U25/U1/clr ) );
    inv_2 \U1213/U916_1_/U25/U1/Ui  ( .x(\y[1] ), .a(\U1213/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_2_/U25/U1/Uclr  ( .x(\U1213/U916_2_/U25/U1/clr ), .a(
        nya), .b(\b[2] ), .c(\d[2] ), .d(\y[2] ) );
    oaoi211_1 \U1213/U916_2_/U25/U1/Uaoi  ( .x(\U1213/U916_2_/U25/U1/ob ), .a(
        \b[2] ), .b(\d[2] ), .c(nya), .d(\U1213/U916_2_/U25/U1/clr ) );
    inv_2 \U1213/U916_2_/U25/U1/Ui  ( .x(\y[2] ), .a(\U1213/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_3_/U25/U1/Uclr  ( .x(\U1213/U916_3_/U25/U1/clr ), .a(
        nya), .b(\b[3] ), .c(\d[3] ), .d(\y[3] ) );
    oaoi211_1 \U1213/U916_3_/U25/U1/Uaoi  ( .x(\U1213/U916_3_/U25/U1/ob ), .a(
        \b[3] ), .b(\d[3] ), .c(nya), .d(\U1213/U916_3_/U25/U1/clr ) );
    inv_2 \U1213/U916_3_/U25/U1/Ui  ( .x(\y[3] ), .a(\U1213/U916_3_/U25/U1/ob 
        ) );
    and3_2 \U1210/U1138/U9  ( .x(\d[3] ), .a(\cdh[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1137/U9  ( .x(\d[2] ), .a(\cdl[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1139/U9  ( .x(\d[1] ), .a(\cdh[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1210/U1136/U9  ( .x(\d[0] ), .a(\cdl[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1162/U1138/U9  ( .x(\a[3] ), .a(ih[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1137/U9  ( .x(\a[2] ), .a(il[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1139/U9  ( .x(\a[1] ), .a(ih[6]), .b(naa), .c(il[7]) );
    and3_2 \U1162/U1136/U9  ( .x(\a[0] ), .a(il[6]), .b(naa), .c(il[7]) );
    and3_2 \U1211/U1138/U9  ( .x(\b[3] ), .a(ih[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1137/U9  ( .x(\b[2] ), .a(il[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1139/U9  ( .x(\b[1] ), .a(ih[4]), .b(nba), .c(il[5]) );
    and3_2 \U1211/U1136/U9  ( .x(\b[0] ), .a(il[4]), .b(nba), .c(il[5]) );
    and3_2 \U1163/U1138/U9  ( .x(\c[3] ), .a(\cdh[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1137/U9  ( .x(\c[2] ), .a(\cdl[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1139/U9  ( .x(\c[1] ), .a(\cdh[2] ), .b(nca), .c(\cdl[3] )
         );
    and3_2 \U1163/U1136/U9  ( .x(\c[0] ), .a(\cdl[2] ), .b(nca), .c(\cdl[3] )
         );
    and2_1 \U1296/U1385/U8  ( .x(cg), .a(nbReset), .b(\U1296/ng ) );
    aoi222_1 \U1296/U1384/U30/U1  ( .x(\U1296/ng ), .a(nca), .b(net195), .c(
        nca), .d(\U1296/U1384/Z ), .e(net195), .f(\U1296/U1384/Z ) );
    inv_1 \U1296/U1384/U30/Uinv  ( .x(\U1296/U1384/Z ), .a(\U1296/ng ) );
    oa31_1 \U1296/U1386/U25/U1/Uclr  ( .x(\U1296/U1386/U25/U1/clr ), .a(
        \twobitack[2] ), .b(cg), .c(nca), .d(net195) );
    oaoi211_1 \U1296/U1386/U25/U1/Uaoi  ( .x(\U1296/U1386/U25/U1/ob ), .a(cg), 
        .b(nca), .c(\twobitack[2] ), .d(\U1296/U1386/U25/U1/clr ) );
    inv_2 \U1296/U1386/U25/U1/Ui  ( .x(net195), .a(\U1296/U1386/U25/U1/ob ) );
    and2_1 \U1298/U1385/U8  ( .x(dg), .a(nbReset), .b(\U1298/ng ) );
    aoi222_1 \U1298/U1384/U30/U1  ( .x(\U1298/ng ), .a(nda), .b(net193), .c(
        nda), .d(\U1298/U1384/Z ), .e(net193), .f(\U1298/U1384/Z ) );
    inv_1 \U1298/U1384/U30/Uinv  ( .x(\U1298/U1384/Z ), .a(\U1298/ng ) );
    oa31_1 \U1298/U1386/U25/U1/Uclr  ( .x(\U1298/U1386/U25/U1/clr ), .a(
        \twobitack[0] ), .b(dg), .c(nda), .d(net193) );
    oaoi211_1 \U1298/U1386/U25/U1/Uaoi  ( .x(\U1298/U1386/U25/U1/ob ), .a(dg), 
        .b(nda), .c(\twobitack[0] ), .d(\U1298/U1386/U25/U1/clr ) );
    inv_2 \U1298/U1386/U25/U1/Ui  ( .x(net193), .a(\U1298/U1386/U25/U1/ob ) );
    and2_1 \U1306/U1385/U8  ( .x(bg), .a(nbReset), .b(\U1306/ng ) );
    aoi222_1 \U1306/U1384/U30/U1  ( .x(\U1306/ng ), .a(nba), .b(\twobitack[1] 
        ), .c(nba), .d(\U1306/U1384/Z ), .e(\twobitack[1] ), .f(
        \U1306/U1384/Z ) );
    inv_1 \U1306/U1384/U30/Uinv  ( .x(\U1306/U1384/Z ), .a(\U1306/ng ) );
    oa31_1 \U1306/U1386/U25/U1/Uclr  ( .x(\U1306/U1386/U25/U1/clr ), .a(net199
        ), .b(bg), .c(nba), .d(\twobitack[1] ) );
    oaoi211_1 \U1306/U1386/U25/U1/Uaoi  ( .x(\U1306/U1386/U25/U1/ob ), .a(bg), 
        .b(nba), .c(net199), .d(\U1306/U1386/U25/U1/clr ) );
    inv_2 \U1306/U1386/U25/U1/Ui  ( .x(\twobitack[1] ), .a(
        \U1306/U1386/U25/U1/ob ) );
    and2_1 \U1295/U1385/U8  ( .x(ag), .a(nbReset), .b(\U1295/ng ) );
    aoi222_1 \U1295/U1384/U30/U1  ( .x(\U1295/ng ), .a(naa), .b(\twobitack[3] 
        ), .c(naa), .d(\U1295/U1384/Z ), .e(\twobitack[3] ), .f(
        \U1295/U1384/Z ) );
    inv_1 \U1295/U1384/U30/Uinv  ( .x(\U1295/U1384/Z ), .a(\U1295/ng ) );
    oa31_1 \U1295/U1386/U25/U1/Uclr  ( .x(\U1295/U1386/U25/U1/clr ), .a(net194
        ), .b(ag), .c(naa), .d(\twobitack[3] ) );
    oaoi211_1 \U1295/U1386/U25/U1/Uaoi  ( .x(\U1295/U1386/U25/U1/ob ), .a(ag), 
        .b(naa), .c(net194), .d(\U1295/U1386/U25/U1/clr ) );
    inv_2 \U1295/U1386/U25/U1/Ui  ( .x(\twobitack[3] ), .a(
        \U1295/U1386/U25/U1/ob ) );
    nand2_1 \U1297/U1131/U5  ( .x(\U1297/s ), .a(\U1297/r ), .b(\U1297/nback )
         );
    nand2_1 \U1297/U1103/U5  ( .x(\U1297/r ), .a(\U1297/naack ), .b(\U1297/s )
         );
    inv_1 \U1297/U1111/U3  ( .x(\U1297/reset ), .a(nbReset) );
    inv_1 \U1297/U1112/U3  ( .x(\U1297/naack ), .a(naa) );
    nor2_1 \U1297/U1130/U5  ( .x(\U1297/nback ), .a(nca), .b(\U1297/reset ) );
    aoai211_1 \U1297/U1128/U28/U1/U1  ( .x(\U1297/U1128/U28/U1/clr ), .a(
        \U1297/r ), .b(\U1297/naack ), .c(cg), .d(csel) );
    nand3_1 \U1297/U1128/U28/U1/U2  ( .x(\U1297/U1128/U28/U1/set ), .a(cg), 
        .b(\U1297/r ), .c(\U1297/naack ) );
    nand2_2 \U1297/U1128/U28/U1/U3  ( .x(csel), .a(\U1297/U1128/U28/U1/clr ), 
        .b(\U1297/U1128/U28/U1/set ) );
    aoai211_1 \U1297/U1127/U28/U1/U1  ( .x(\U1297/U1127/U28/U1/clr ), .a(
        \U1297/s ), .b(\U1297/nback ), .c(ag), .d(asel) );
    nand3_1 \U1297/U1127/U28/U1/U2  ( .x(\U1297/U1127/U28/U1/set ), .a(ag), 
        .b(\U1297/s ), .c(\U1297/nback ) );
    nand2_2 \U1297/U1127/U28/U1/U3  ( .x(asel), .a(\U1297/U1127/U28/U1/clr ), 
        .b(\U1297/U1127/U28/U1/set ) );
    nand2_1 \U1300/U1131/U5  ( .x(\U1300/s ), .a(\U1300/r ), .b(\U1300/nback )
         );
    nand2_1 \U1300/U1103/U5  ( .x(\U1300/r ), .a(\U1300/naack ), .b(\U1300/s )
         );
    inv_1 \U1300/U1111/U3  ( .x(\U1300/reset ), .a(nbReset) );
    inv_1 \U1300/U1112/U3  ( .x(\U1300/naack ), .a(nba) );
    nor2_1 \U1300/U1130/U5  ( .x(\U1300/nback ), .a(nda), .b(\U1300/reset ) );
    aoai211_1 \U1300/U1128/U28/U1/U1  ( .x(\U1300/U1128/U28/U1/clr ), .a(
        \U1300/r ), .b(\U1300/naack ), .c(dg), .d(dsel) );
    nand3_1 \U1300/U1128/U28/U1/U2  ( .x(\U1300/U1128/U28/U1/set ), .a(dg), 
        .b(\U1300/r ), .c(\U1300/naack ) );
    nand2_2 \U1300/U1128/U28/U1/U3  ( .x(dsel), .a(\U1300/U1128/U28/U1/clr ), 
        .b(\U1300/U1128/U28/U1/set ) );
    aoai211_1 \U1300/U1127/U28/U1/U1  ( .x(\U1300/U1127/U28/U1/clr ), .a(
        \U1300/s ), .b(\U1300/nback ), .c(bg), .d(bsel) );
    nand3_1 \U1300/U1127/U28/U1/U2  ( .x(\U1300/U1127/U28/U1/set ), .a(bg), 
        .b(\U1300/s ), .c(\U1300/nback ) );
    nand2_2 \U1300/U1127/U28/U1/U3  ( .x(bsel), .a(\U1300/U1127/U28/U1/clr ), 
        .b(\U1300/U1127/U28/U1/set ) );
    aoai211_1 \U1289/U1150/U28/U1/U1  ( .x(\U1289/U1150/U28/U1/clr ), .a(il[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[2] ) );
    nand3_1 \U1289/U1150/U28/U1/U2  ( .x(\U1289/U1150/U28/U1/set ), .a(net195), 
        .b(il[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1150/U28/U1/U3  ( .x(\cdl[2] ), .a(
        \U1289/U1150/U28/U1/clr ), .b(\U1289/U1150/U28/U1/set ) );
    aoai211_1 \U1289/U1152/U28/U1/U1  ( .x(\U1289/U1152/U28/U1/clr ), .a(il[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[3] ) );
    nand3_1 \U1289/U1152/U28/U1/U2  ( .x(\U1289/U1152/U28/U1/set ), .a(net195), 
        .b(il[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1152/U28/U1/U3  ( .x(\cdl[3] ), .a(
        \U1289/U1152/U28/U1/clr ), .b(\U1289/U1152/U28/U1/set ) );
    aoai211_1 \U1289/U1149/U28/U1/U1  ( .x(\U1289/U1149/U28/U1/clr ), .a(ih[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[2] ) );
    nand3_1 \U1289/U1149/U28/U1/U2  ( .x(\U1289/U1149/U28/U1/set ), .a(net195), 
        .b(ih[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1149/U28/U1/U3  ( .x(\cdh[2] ), .a(
        \U1289/U1149/U28/U1/clr ), .b(\U1289/U1149/U28/U1/set ) );
    aoai211_1 \U1289/U1151/U28/U1/U1  ( .x(\U1289/U1151/U28/U1/clr ), .a(ih[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[3] ) );
    nand3_1 \U1289/U1151/U28/U1/U2  ( .x(\U1289/U1151/U28/U1/set ), .a(net195), 
        .b(ih[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1151/U28/U1/U3  ( .x(\cdh[3] ), .a(
        \U1289/U1151/U28/U1/clr ), .b(\U1289/U1151/U28/U1/set ) );
    inv_1 \U1289/U1148/U1147/U3  ( .x(\U1289/U1148/net189 ), .a(
        \U1289/bnreset ) );
    nor2_1 \U1289/U1148/U582/U5  ( .x(\U1289/U1148/net192 ), .a(\cdl[3] ), .b(
        \cdh[3] ) );
    nor2_1 \U1289/U1148/U580/U5  ( .x(\U1289/U1148/net191 ), .a(\cdl[2] ), .b(
        \cdh[2] ) );
    nor2_2 \U1289/U1148/U1146/U6  ( .x(\twobitack[2] ), .a(
        \U1289/U1148/net190 ), .b(\U1289/U1148/net189 ) );
    aoi222_1 \U1289/U1148/U1141/U30/U1  ( .x(\U1289/U1148/net190 ), .a(
        \U1289/U1148/net191 ), .b(\U1289/U1148/net192 ), .c(
        \U1289/U1148/net191 ), .d(\U1289/U1148/U1141/Z ), .e(
        \U1289/U1148/net192 ), .f(\U1289/U1148/U1141/Z ) );
    inv_1 \U1289/U1148/U1141/U30/Uinv  ( .x(\U1289/U1148/U1141/Z ), .a(
        \U1289/U1148/net190 ) );
    aoai211_1 \U1271/U1150/U28/U1/U1  ( .x(\U1271/U1150/U28/U1/clr ), .a(il[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[0] ) );
    nand3_1 \U1271/U1150/U28/U1/U2  ( .x(\U1271/U1150/U28/U1/set ), .a(net193), 
        .b(il[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1150/U28/U1/U3  ( .x(\cdl[0] ), .a(
        \U1271/U1150/U28/U1/clr ), .b(\U1271/U1150/U28/U1/set ) );
    aoai211_1 \U1271/U1152/U28/U1/U1  ( .x(\U1271/U1152/U28/U1/clr ), .a(il[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[1] ) );
    nand3_1 \U1271/U1152/U28/U1/U2  ( .x(\U1271/U1152/U28/U1/set ), .a(net193), 
        .b(il[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1152/U28/U1/U3  ( .x(\cdl[1] ), .a(
        \U1271/U1152/U28/U1/clr ), .b(\U1271/U1152/U28/U1/set ) );
    aoai211_1 \U1271/U1149/U28/U1/U1  ( .x(\U1271/U1149/U28/U1/clr ), .a(ih[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[0] ) );
    nand3_1 \U1271/U1149/U28/U1/U2  ( .x(\U1271/U1149/U28/U1/set ), .a(net193), 
        .b(ih[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1149/U28/U1/U3  ( .x(\cdh[0] ), .a(
        \U1271/U1149/U28/U1/clr ), .b(\U1271/U1149/U28/U1/set ) );
    aoai211_1 \U1271/U1151/U28/U1/U1  ( .x(\U1271/U1151/U28/U1/clr ), .a(ih[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[1] ) );
    nand3_1 \U1271/U1151/U28/U1/U2  ( .x(\U1271/U1151/U28/U1/set ), .a(net193), 
        .b(ih[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1151/U28/U1/U3  ( .x(\cdh[1] ), .a(
        \U1271/U1151/U28/U1/clr ), .b(\U1271/U1151/U28/U1/set ) );
    inv_1 \U1271/U1148/U1147/U3  ( .x(\U1271/U1148/net189 ), .a(
        \U1271/bnreset ) );
    nor2_1 \U1271/U1148/U582/U5  ( .x(\U1271/U1148/net192 ), .a(\cdl[1] ), .b(
        \cdh[1] ) );
    nor2_1 \U1271/U1148/U580/U5  ( .x(\U1271/U1148/net191 ), .a(\cdl[0] ), .b(
        \cdh[0] ) );
    nor2_2 \U1271/U1148/U1146/U6  ( .x(\twobitack[0] ), .a(
        \U1271/U1148/net190 ), .b(\U1271/U1148/net189 ) );
    aoi222_1 \U1271/U1148/U1141/U30/U1  ( .x(\U1271/U1148/net190 ), .a(
        \U1271/U1148/net191 ), .b(\U1271/U1148/net192 ), .c(
        \U1271/U1148/net191 ), .d(\U1271/U1148/U1141/Z ), .e(
        \U1271/U1148/net192 ), .f(\U1271/U1148/U1141/Z ) );
    inv_1 \U1271/U1148/U1141/U30/Uinv  ( .x(\U1271/U1148/U1141/Z ), .a(
        \U1271/U1148/net190 ) );
    nand2_1 \U1225/U1128/U5  ( .x(\U1225/s ), .a(\U1225/r ), .b(\U1225/nback )
         );
    nand2_1 \U1225/U1103/U5  ( .x(\U1225/r ), .a(\U1225/naack ), .b(\U1225/s )
         );
    inv_1 \U1225/U1111/U3  ( .x(\U1225/reset ), .a(nbReset) );
    inv_1 \U1225/U1112/U3  ( .x(\U1225/naack ), .a(nxa) );
    nor2_1 \U1225/U1127/U5  ( .x(\U1225/nback ), .a(nyla), .b(\U1225/reset )
         );
    and2_2 \U1225/U1129/U8  ( .x(xsel), .a(\U1225/nback ), .b(\U1225/s ) );
    and2_2 \U1225/U1124/U8  ( .x(ysel), .a(\U1225/r ), .b(\U1225/naack ) );
    and3_4 \U1308/U20/U9  ( .x(nya), .a(\U1308/nack[1] ), .b(\U1308/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U1308/U18/U5  ( .x(\U1308/nack[0] ), .a(\yl[3] ), .b(\yl[0] ) );
    nor2_1 \U1308/U19/U5  ( .x(\U1308/nack[1] ), .a(\yl[1] ), .b(\yl[2] ) );
    ao222_2 \U1308/U15_0_/U19/U1/U1  ( .x(\yl[0] ), .a(\y[0] ), .b(nyla), .c(
        \y[0] ), .d(\yl[0] ), .e(nyla), .f(\yl[0] ) );
    ao222_2 \U1308/U15_1_/U19/U1/U1  ( .x(\yl[1] ), .a(\y[1] ), .b(nyla), .c(
        \y[1] ), .d(\yl[1] ), .e(nyla), .f(\yl[1] ) );
    ao222_2 \U1308/U15_2_/U19/U1/U1  ( .x(\yl[2] ), .a(\y[2] ), .b(nyla), .c(
        \y[2] ), .d(\yl[2] ), .e(nyla), .f(\yl[2] ) );
    ao222_2 \U1308/U15_3_/U19/U1/U1  ( .x(\yl[3] ), .a(\y[3] ), .b(nyla), .c(
        \y[3] ), .d(\yl[3] ), .e(nyla), .f(\yl[3] ) );
    buf_3 U1 ( .x(\U1271/bnreset ), .a(nbReset) );
    buf_3 U2 ( .x(\U1289/bnreset ), .a(nbReset) );
endmodule


module chain_mergepackets_1 ( naa, nba, o, a, b, nReset, noa );
output [4:0] o;
input  [4:0] a;
input  [4:0] b;
input  nReset, noa;
output naa, nba;
    wire \noack[1] , \noack[0] , reset, bsel, as, setb, asel, seta, 
        \U916_0_/U25/U1/clr , \U916_0_/U25/U1/ob , \U916_1_/U25/U1/clr , 
        \U916_1_/U25/U1/ob , \U916_2_/U25/U1/clr , \U916_2_/U25/U1/ob , 
        \U916_3_/U25/U1/clr , \U916_3_/U25/U1/ob ;
    and2_1 \U1155/U8  ( .x(as), .a(seta), .b(asel) );
    nand2_1 \U1145/U5  ( .x(asel), .a(bsel), .b(seta) );
    nand2_1 \U1103/U5  ( .x(bsel), .a(setb), .b(asel) );
    inv_1 \U1135/U3  ( .x(reset), .a(nReset) );
    inv_1 \U1134/U3  ( .x(setb), .a(a[4]) );
    and3_2 \U1154/U9  ( .x(naa), .a(\noack[1] ), .b(\noack[0] ), .c(as) );
    nor3_1 \U1127/U7  ( .x(\noack[0] ), .a(o[1]), .b(reset), .c(o[0]) );
    nor2_1 \U1132/U5  ( .x(\noack[1] ), .a(o[3]), .b(o[2]) );
    oa31_1 \U916_0_/U25/U1/Uclr  ( .x(\U916_0_/U25/U1/clr ), .a(noa), .b(a[0]), 
        .c(b[0]), .d(o[0]) );
    oaoi211_1 \U916_0_/U25/U1/Uaoi  ( .x(\U916_0_/U25/U1/ob ), .a(a[0]), .b(b
        [0]), .c(noa), .d(\U916_0_/U25/U1/clr ) );
    inv_2 \U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U916_0_/U25/U1/ob ) );
    oa31_1 \U916_1_/U25/U1/Uclr  ( .x(\U916_1_/U25/U1/clr ), .a(noa), .b(a[1]), 
        .c(b[1]), .d(o[1]) );
    oaoi211_1 \U916_1_/U25/U1/Uaoi  ( .x(\U916_1_/U25/U1/ob ), .a(a[1]), .b(b
        [1]), .c(noa), .d(\U916_1_/U25/U1/clr ) );
    inv_2 \U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U916_1_/U25/U1/ob ) );
    oa31_1 \U916_2_/U25/U1/Uclr  ( .x(\U916_2_/U25/U1/clr ), .a(noa), .b(a[2]), 
        .c(b[2]), .d(o[2]) );
    oaoi211_1 \U916_2_/U25/U1/Uaoi  ( .x(\U916_2_/U25/U1/ob ), .a(a[2]), .b(b
        [2]), .c(noa), .d(\U916_2_/U25/U1/clr ) );
    inv_2 \U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U916_2_/U25/U1/ob ) );
    oa31_1 \U916_3_/U25/U1/Uclr  ( .x(\U916_3_/U25/U1/clr ), .a(noa), .b(a[3]), 
        .c(b[3]), .d(o[3]) );
    oaoi211_1 \U916_3_/U25/U1/Uaoi  ( .x(\U916_3_/U25/U1/ob ), .a(a[3]), .b(b
        [3]), .c(noa), .d(\U916_3_/U25/U1/clr ) );
    inv_2 \U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U916_3_/U25/U1/ob ) );
    ao222_2 \U1148/U19/U1/U1  ( .x(o[4]), .a(noa), .b(b[4]), .c(noa), .d(o[4]), 
        .e(b[4]), .f(o[4]) );
    aoi21_1 \U1153/U11  ( .x(seta), .a(o[4]), .b(setb), .c(reset) );
    and3_3 U1 ( .x(nba), .a(bsel), .b(\noack[0] ), .c(\noack[1] ) );
endmodule


module initiator_dport ( cack, chaincommand, err, nchainresponseack, nrouteack, 
    rd, routetxreq, rrnw, a, chainresponse, col, crnw, itag, lock, nReset, 
    nchaincommandack, pred, rack, route, routetxack, seq, size, wd );
output [4:0] chaincommand;
output [1:0] err;
output [63:0] rd;
output [1:0] rrnw;
input  [63:0] a;
input  [4:0] chainresponse;
input  [5:0] col;
input  [1:0] crnw;
input  [9:0] itag;
input  [1:0] lock;
input  [1:0] pred;
input  [4:0] route;
input  [1:0] seq;
input  [3:0] size;
input  [63:0] wd;
input  nReset, nchaincommandack, rack, routetxack;
output cack, nchainresponseack, nrouteack, routetxreq;
    wire \irbh[7] , \irbh[6] , \irbh[5] , \irbh[4] , \irbh[3] , \irbh[2] , 
        \irbh[1] , \irbh[0] , \ipayload[4] , \ipayload[3] , \ipayload[2] , 
        \ipayload[1] , \ipayload[0] , \icbh[7] , \icbh[6] , \icbh[5] , 
        \icbh[4] , \icbh[3] , \icbh[2] , \icbh[1] , \icbh[0] , \cstatus[1] , 
        \cstatus[0] , \irbl[7] , \irbl[6] , \irbl[5] , \irbl[4] , \irbl[3] , 
        \irbl[2] , \irbl[1] , \irbl[0] , \rstatus[1] , \rstatus[0] , 
        \can_defer[0] , \icbl[7] , \icbl[6] , \icbl[5] , \icbl[4] , \icbl[3] , 
        \icbl[2] , \icbl[1] , \icbl[0] , nircba, nResetb, responseack, 
        rstatusack, net165, reset, tok_ack, net170, ictrlack, icmdack, 
        ncstatusack, net116, pltxreq, net115, net128, pltxack, nicba, 
        nipayloadack, \U1662/U28/U1/clr , \U1662/U28/U1/set ;
    chain_irdemuxNew_1 U1442 ( .err(err), .ncback(nircba), .rd(rd), .rnw(rrnw), 
        .status({\rstatus[1] , \rstatus[0] }), .cbh({\irbh[7] , \irbh[6] , 
        \irbh[5] , \irbh[4] , \irbh[3] , \irbh[2] , \irbh[1] , \irbh[0] }), 
        .cbl({\irbl[7] , \irbl[6] , \irbl[5] , \irbl[4] , \irbl[3] , \irbl[2] , 
        \irbl[1] , \irbl[0] }), .nReset(nResetb), .nack(responseack), 
        .statusack(rstatusack) );
    chain_fr2dr_byte_4 chain_decoder ( .nia(nchainresponseack), .oh({\irbh[7] , 
        \irbh[6] , \irbh[5] , \irbh[4] , \irbh[3] , \irbh[2] , \irbh[1] , 
        \irbh[0] }), .ol({\irbl[7] , \irbl[6] , \irbl[5] , \irbl[4] , 
        \irbl[3] , \irbl[2] , \irbl[1] , \irbl[0] }), .i(chainresponse), 
        .nReset(nResetb), .noa(nircba) );
    chain_ic_ctrl_1 cmd_ctrl ( .ack(ictrlack), .candefer(\can_defer[0] ), 
        .eop(net116), .nstatack(ncstatusack), .pltxreq(pltxreq), .routetxreq(
        routetxreq), .tok_ack(tok_ack), .accept(\cstatus[0] ), .candefer_ack({
        1'b0, \can_defer[0] }), .defer(\cstatus[1] ), .eopack(net115), .lock(
        lock), .nReset(net128), .pltxack(pltxack), .routetxack(routetxack), 
        .tok_err(err[1]), .tok_ok(err[0]) );
    chain_icmux_1 cmd_mux ( .ack(icmdack), .chainh({\icbh[7] , \icbh[6] , 
        \icbh[5] , \icbh[4] , \icbh[3] , \icbh[2] , \icbh[1] , \icbh[0] }), 
        .chainl({\icbl[7] , \icbl[6] , \icbl[5] , \icbl[4] , \icbl[3] , 
        \icbl[2] , \icbl[1] , \icbl[0] }), .sendack(pltxack), .addr(a), .col(
        col), .itag(itag), .lock(lock), .nReset(net128), .nia(nicba), .pred(
        pred), .rnw(crnw), .sendreq(pltxreq), .seq(seq), .size(size), .wd(wd)
         );
    chain_dr2fr_byte_1 U1604 ( .eop_ack(net115), .ia(nicba), .o({\ipayload[4] , 
        \ipayload[3] , \ipayload[2] , \ipayload[1] , \ipayload[0] }), .eop(
        net116), .ih({\icbh[7] , \icbh[6] , \icbh[5] , \icbh[4] , \icbh[3] , 
        \icbh[2] , \icbh[1] , \icbh[0] }), .il({\icbl[7] , \icbl[6] , 
        \icbl[5] , \icbl[4] , \icbl[3] , \icbl[2] , \icbl[1] , \icbl[0] }), 
        .nReset(net128), .noa(nipayloadack) );
    chain_mergepackets_1 U1605 ( .naa(nrouteack), .nba(nipayloadack), .o(
        chaincommand), .a(route), .b({\ipayload[4] , \ipayload[3] , 
        \ipayload[2] , \ipayload[1] , \ipayload[0] }), .nReset(net128), .noa(
        nchaincommandack) );
    and2_1 U1676 ( .x(cack), .a(net170), .b(nResetb) );
    inv_4 \U1643/U3  ( .x(net128), .a(reset) );
    or2_4 \U1660/U12  ( .x(net165), .a(\cstatus[0] ), .b(\cstatus[1] ) );
    or2_1 \U1661/U12  ( .x(rstatusack), .a(net165), .b(reset) );
    ao222_2 \status_pipe_0_/U19/U1/U1  ( .x(\cstatus[0] ), .a(\rstatus[0] ), 
        .b(ncstatusack), .c(\rstatus[0] ), .d(\cstatus[0] ), .e(ncstatusack), 
        .f(\cstatus[0] ) );
    ao222_2 \status_pipe_1_/U19/U1/U1  ( .x(\cstatus[1] ), .a(\rstatus[1] ), 
        .b(ncstatusack), .c(\rstatus[1] ), .d(\cstatus[1] ), .e(ncstatusack), 
        .f(\cstatus[1] ) );
    ao222_1 \U1609/U18/U1/U1  ( .x(net170), .a(ictrlack), .b(icmdack), .c(
        ictrlack), .d(net170), .e(icmdack), .f(net170) );
    aoai211_1 \U1662/U28/U1/U1  ( .x(\U1662/U28/U1/clr ), .a(rack), .b(nResetb
        ), .c(tok_ack), .d(responseack) );
    nand3_1 \U1662/U28/U1/U2  ( .x(\U1662/U28/U1/set ), .a(tok_ack), .b(rack), 
        .c(nResetb) );
    nand2_2 \U1662/U28/U1/U3  ( .x(responseack), .a(\U1662/U28/U1/clr ), .b(
        \U1662/U28/U1/set ) );
    inv_2 U1 ( .x(reset), .a(nResetb) );
    buf_3 U2 ( .x(nResetb), .a(nReset) );
endmodule


module matched_delay_m2cp_com_dport ( x, a );
input  a;
output x;
    wire n2;
    buf_1 I1 ( .x(n2), .a(a) );
    buf_16 U1 ( .x(x), .a(n2) );
endmodule


module matched_delay_m2cp_resp_dport ( x, a );
input  a;
output x;
    assign x = a;
endmodule


module sr2dr_word_2 ( i, req, h, l );
input  [31:0] i;
output [31:0] h;
output [31:0] l;
input  req;
    wire \U31/nl , \U31/ni , \U31/nh , \U30/nl , \U30/ni , \U30/nh , \U29/nl , 
        \U29/ni , \U29/nh , \U28/nl , \U28/ni , \U28/nh , \U27/nl , \U27/ni , 
        \U27/nh , \U26/nl , \U26/ni , \U26/nh , \U25/nl , \U25/ni , \U25/nh , 
        \U24/nl , \U24/ni , \U24/nh , \U23/nl , \U23/ni , \U23/nh , \U22/nl , 
        \U22/ni , \U22/nh , \U21/nl , \U21/ni , \U21/nh , \U20/nl , \U20/ni , 
        \U20/nh , \U19/nl , \U19/ni , \U19/nh , \U18/nl , \U18/ni , \U18/nh , 
        \U17/nl , \U17/ni , \U17/nh , \U16/nl , \U16/ni , \U16/nh , \U15/nl , 
        \U15/ni , \U15/nh , \U14/nl , \U14/ni , \U14/nh , \U13/nl , \U13/ni , 
        \U13/nh , \U12/nl , \U12/ni , \U12/nh , \U11/nl , \U11/ni , \U11/nh , 
        \U10/nl , \U10/ni , \U10/nh , \U9/nl , \U9/ni , \U9/nh , \U8/nl , 
        \U8/ni , \U8/nh , \U7/nl , \U7/ni , \U7/nh , \U6/nl , \U6/ni , \U6/nh , 
        \U5/nl , \U5/ni , \U5/nh , \U4/nl , \U4/ni , \U4/nh , \U3/nl , \U3/ni , 
        \U3/nh , \U2/nl , \U2/ni , \U2/nh , \U1/nl , \U1/ni , \U1/nh , \U0/nl , 
        \U0/ni , \U0/nh , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
    inv_1 \U31/Uii  ( .x(\U31/ni ), .a(i[31]) );
    inv_1 \U31/Uih  ( .x(\U31/nh ), .a(h[31]) );
    inv_1 \U31/Uil  ( .x(\U31/nl ), .a(l[31]) );
    ao23_1 \U31/Ucl/U1/U1  ( .x(l[31]), .a(n9), .b(l[31]), .c(n1), .d(\U31/ni 
        ), .e(\U31/nh ) );
    ao23_1 \U31/Uch/U1/U1  ( .x(h[31]), .a(n9), .b(h[31]), .c(n2), .d(i[31]), 
        .e(\U31/nl ) );
    inv_1 \U30/Uii  ( .x(\U30/ni ), .a(i[30]) );
    inv_1 \U30/Uih  ( .x(\U30/nh ), .a(h[30]) );
    inv_1 \U30/Uil  ( .x(\U30/nl ), .a(l[30]) );
    ao23_1 \U30/Ucl/U1/U1  ( .x(l[30]), .a(n8), .b(l[30]), .c(n1), .d(\U30/ni 
        ), .e(\U30/nh ) );
    ao23_1 \U30/Uch/U1/U1  ( .x(h[30]), .a(n8), .b(h[30]), .c(n1), .d(i[30]), 
        .e(\U30/nl ) );
    inv_1 \U29/Uii  ( .x(\U29/ni ), .a(i[29]) );
    inv_1 \U29/Uih  ( .x(\U29/nh ), .a(h[29]) );
    inv_1 \U29/Uil  ( .x(\U29/nl ), .a(l[29]) );
    ao23_1 \U29/Ucl/U1/U1  ( .x(l[29]), .a(n8), .b(l[29]), .c(n1), .d(\U29/ni 
        ), .e(\U29/nh ) );
    ao23_1 \U29/Uch/U1/U1  ( .x(h[29]), .a(n8), .b(h[29]), .c(n2), .d(i[29]), 
        .e(\U29/nl ) );
    inv_1 \U28/Uii  ( .x(\U28/ni ), .a(i[28]) );
    inv_1 \U28/Uih  ( .x(\U28/nh ), .a(h[28]) );
    inv_1 \U28/Uil  ( .x(\U28/nl ), .a(l[28]) );
    ao23_1 \U28/Ucl/U1/U1  ( .x(l[28]), .a(n8), .b(l[28]), .c(n2), .d(\U28/ni 
        ), .e(\U28/nh ) );
    ao23_1 \U28/Uch/U1/U1  ( .x(h[28]), .a(n8), .b(h[28]), .c(n2), .d(i[28]), 
        .e(\U28/nl ) );
    inv_1 \U27/Uii  ( .x(\U27/ni ), .a(i[27]) );
    inv_1 \U27/Uih  ( .x(\U27/nh ), .a(h[27]) );
    inv_1 \U27/Uil  ( .x(\U27/nl ), .a(l[27]) );
    ao23_1 \U27/Ucl/U1/U1  ( .x(l[27]), .a(n8), .b(l[27]), .c(n2), .d(\U27/ni 
        ), .e(\U27/nh ) );
    ao23_1 \U27/Uch/U1/U1  ( .x(h[27]), .a(n8), .b(h[27]), .c(n2), .d(i[27]), 
        .e(\U27/nl ) );
    inv_1 \U26/Uii  ( .x(\U26/ni ), .a(i[26]) );
    inv_1 \U26/Uih  ( .x(\U26/nh ), .a(h[26]) );
    inv_1 \U26/Uil  ( .x(\U26/nl ), .a(l[26]) );
    ao23_1 \U26/Ucl/U1/U1  ( .x(l[26]), .a(n7), .b(l[26]), .c(n2), .d(\U26/ni 
        ), .e(\U26/nh ) );
    ao23_1 \U26/Uch/U1/U1  ( .x(h[26]), .a(n7), .b(h[26]), .c(n4), .d(i[26]), 
        .e(\U26/nl ) );
    inv_1 \U25/Uii  ( .x(\U25/ni ), .a(i[25]) );
    inv_1 \U25/Uih  ( .x(\U25/nh ), .a(h[25]) );
    inv_1 \U25/Uil  ( .x(\U25/nl ), .a(l[25]) );
    ao23_1 \U25/Ucl/U1/U1  ( .x(l[25]), .a(n7), .b(l[25]), .c(n4), .d(\U25/ni 
        ), .e(\U25/nh ) );
    ao23_1 \U25/Uch/U1/U1  ( .x(h[25]), .a(n7), .b(h[25]), .c(n4), .d(i[25]), 
        .e(\U25/nl ) );
    inv_1 \U24/Uii  ( .x(\U24/ni ), .a(i[24]) );
    inv_1 \U24/Uih  ( .x(\U24/nh ), .a(h[24]) );
    inv_1 \U24/Uil  ( .x(\U24/nl ), .a(l[24]) );
    ao23_1 \U24/Ucl/U1/U1  ( .x(l[24]), .a(n7), .b(l[24]), .c(n4), .d(\U24/ni 
        ), .e(\U24/nh ) );
    ao23_1 \U24/Uch/U1/U1  ( .x(h[24]), .a(n7), .b(h[24]), .c(n4), .d(i[24]), 
        .e(\U24/nl ) );
    inv_1 \U23/Uii  ( .x(\U23/ni ), .a(i[23]) );
    inv_1 \U23/Uih  ( .x(\U23/nh ), .a(h[23]) );
    inv_1 \U23/Uil  ( .x(\U23/nl ), .a(l[23]) );
    ao23_1 \U23/Ucl/U1/U1  ( .x(l[23]), .a(n7), .b(l[23]), .c(n3), .d(\U23/ni 
        ), .e(\U23/nh ) );
    ao23_1 \U23/Uch/U1/U1  ( .x(h[23]), .a(n7), .b(h[23]), .c(n3), .d(i[23]), 
        .e(\U23/nl ) );
    inv_1 \U22/Uii  ( .x(\U22/ni ), .a(i[22]) );
    inv_1 \U22/Uih  ( .x(\U22/nh ), .a(h[22]) );
    inv_1 \U22/Uil  ( .x(\U22/nl ), .a(l[22]) );
    ao23_1 \U22/Ucl/U1/U1  ( .x(l[22]), .a(n6), .b(l[22]), .c(n3), .d(\U22/ni 
        ), .e(\U22/nh ) );
    ao23_1 \U22/Uch/U1/U1  ( .x(h[22]), .a(n6), .b(h[22]), .c(n3), .d(i[22]), 
        .e(\U22/nl ) );
    inv_1 \U21/Uii  ( .x(\U21/ni ), .a(i[21]) );
    inv_1 \U21/Uih  ( .x(\U21/nh ), .a(h[21]) );
    inv_1 \U21/Uil  ( .x(\U21/nl ), .a(l[21]) );
    ao23_1 \U21/Ucl/U1/U1  ( .x(l[21]), .a(n6), .b(l[21]), .c(n3), .d(\U21/ni 
        ), .e(\U21/nh ) );
    ao23_1 \U21/Uch/U1/U1  ( .x(h[21]), .a(n6), .b(h[21]), .c(n3), .d(i[21]), 
        .e(\U21/nl ) );
    inv_1 \U20/Uii  ( .x(\U20/ni ), .a(i[20]) );
    inv_1 \U20/Uih  ( .x(\U20/nh ), .a(h[20]) );
    inv_1 \U20/Uil  ( .x(\U20/nl ), .a(l[20]) );
    ao23_1 \U20/Ucl/U1/U1  ( .x(l[20]), .a(n6), .b(l[20]), .c(n5), .d(\U20/ni 
        ), .e(\U20/nh ) );
    ao23_1 \U20/Uch/U1/U1  ( .x(h[20]), .a(n6), .b(h[20]), .c(n4), .d(i[20]), 
        .e(\U20/nl ) );
    inv_1 \U19/Uii  ( .x(\U19/ni ), .a(i[19]) );
    inv_1 \U19/Uih  ( .x(\U19/nh ), .a(h[19]) );
    inv_1 \U19/Uil  ( .x(\U19/nl ), .a(l[19]) );
    ao23_1 \U19/Ucl/U1/U1  ( .x(l[19]), .a(n6), .b(l[19]), .c(n4), .d(\U19/ni 
        ), .e(\U19/nh ) );
    ao23_1 \U19/Uch/U1/U1  ( .x(h[19]), .a(n6), .b(h[19]), .c(n4), .d(i[19]), 
        .e(\U19/nl ) );
    inv_1 \U18/Uii  ( .x(\U18/ni ), .a(i[18]) );
    inv_1 \U18/Uih  ( .x(\U18/nh ), .a(h[18]) );
    inv_1 \U18/Uil  ( .x(\U18/nl ), .a(l[18]) );
    ao23_1 \U18/Ucl/U1/U1  ( .x(l[18]), .a(n5), .b(l[18]), .c(n5), .d(\U18/ni 
        ), .e(\U18/nh ) );
    ao23_1 \U18/Uch/U1/U1  ( .x(h[18]), .a(n5), .b(h[18]), .c(n5), .d(i[18]), 
        .e(\U18/nl ) );
    inv_1 \U17/Uii  ( .x(\U17/ni ), .a(i[17]) );
    inv_1 \U17/Uih  ( .x(\U17/nh ), .a(h[17]) );
    inv_1 \U17/Uil  ( .x(\U17/nl ), .a(l[17]) );
    ao23_1 \U17/Ucl/U1/U1  ( .x(l[17]), .a(n6), .b(l[17]), .c(n5), .d(\U17/ni 
        ), .e(\U17/nh ) );
    ao23_1 \U17/Uch/U1/U1  ( .x(h[17]), .a(n7), .b(h[17]), .c(n4), .d(i[17]), 
        .e(\U17/nl ) );
    inv_1 \U16/Uii  ( .x(\U16/ni ), .a(i[16]) );
    inv_1 \U16/Uih  ( .x(\U16/nh ), .a(h[16]) );
    inv_1 \U16/Uil  ( .x(\U16/nl ), .a(l[16]) );
    ao23_1 \U16/Ucl/U1/U1  ( .x(l[16]), .a(n9), .b(l[16]), .c(n3), .d(\U16/ni 
        ), .e(\U16/nh ) );
    ao23_1 \U16/Uch/U1/U1  ( .x(h[16]), .a(n9), .b(h[16]), .c(n1), .d(i[16]), 
        .e(\U16/nl ) );
    inv_1 \U15/Uii  ( .x(\U15/ni ), .a(i[15]) );
    inv_1 \U15/Uih  ( .x(\U15/nh ), .a(h[15]) );
    inv_1 \U15/Uil  ( .x(\U15/nl ), .a(l[15]) );
    ao23_1 \U15/Ucl/U1/U1  ( .x(l[15]), .a(n8), .b(l[15]), .c(n1), .d(\U15/ni 
        ), .e(\U15/nh ) );
    ao23_1 \U15/Uch/U1/U1  ( .x(h[15]), .a(n7), .b(h[15]), .c(n1), .d(i[15]), 
        .e(\U15/nl ) );
    inv_1 \U14/Uii  ( .x(\U14/ni ), .a(i[14]) );
    inv_1 \U14/Uih  ( .x(\U14/nh ), .a(h[14]) );
    inv_1 \U14/Uil  ( .x(\U14/nl ), .a(l[14]) );
    ao23_1 \U14/Ucl/U1/U1  ( .x(l[14]), .a(n6), .b(l[14]), .c(n1), .d(\U14/ni 
        ), .e(\U14/nh ) );
    ao23_1 \U14/Uch/U1/U1  ( .x(h[14]), .a(n6), .b(h[14]), .c(n3), .d(i[14]), 
        .e(\U14/nl ) );
    inv_1 \U13/Uii  ( .x(\U13/ni ), .a(i[13]) );
    inv_1 \U13/Uih  ( .x(\U13/nh ), .a(h[13]) );
    inv_1 \U13/Uil  ( .x(\U13/nl ), .a(l[13]) );
    ao23_1 \U13/Ucl/U1/U1  ( .x(l[13]), .a(n6), .b(l[13]), .c(n4), .d(\U13/ni 
        ), .e(\U13/nh ) );
    ao23_1 \U13/Uch/U1/U1  ( .x(h[13]), .a(n6), .b(h[13]), .c(n4), .d(i[13]), 
        .e(\U13/nl ) );
    inv_1 \U12/Uii  ( .x(\U12/ni ), .a(i[12]) );
    inv_1 \U12/Uih  ( .x(\U12/nh ), .a(h[12]) );
    inv_1 \U12/Uil  ( .x(\U12/nl ), .a(l[12]) );
    ao23_1 \U12/Ucl/U1/U1  ( .x(l[12]), .a(n5), .b(l[12]), .c(n4), .d(\U12/ni 
        ), .e(\U12/nh ) );
    ao23_1 \U12/Uch/U1/U1  ( .x(h[12]), .a(n5), .b(h[12]), .c(n4), .d(i[12]), 
        .e(\U12/nl ) );
    inv_1 \U11/Uii  ( .x(\U11/ni ), .a(i[11]) );
    inv_1 \U11/Uih  ( .x(\U11/nh ), .a(h[11]) );
    inv_1 \U11/Uil  ( .x(\U11/nl ), .a(l[11]) );
    ao23_1 \U11/Ucl/U1/U1  ( .x(l[11]), .a(n5), .b(l[11]), .c(n4), .d(\U11/ni 
        ), .e(\U11/nh ) );
    ao23_1 \U11/Uch/U1/U1  ( .x(h[11]), .a(n5), .b(h[11]), .c(n4), .d(i[11]), 
        .e(\U11/nl ) );
    inv_1 \U10/Uii  ( .x(\U10/ni ), .a(i[10]) );
    inv_1 \U10/Uih  ( .x(\U10/nh ), .a(h[10]) );
    inv_1 \U10/Uil  ( .x(\U10/nl ), .a(l[10]) );
    ao23_1 \U10/Ucl/U1/U1  ( .x(l[10]), .a(n5), .b(l[10]), .c(n3), .d(\U10/ni 
        ), .e(\U10/nh ) );
    ao23_1 \U10/Uch/U1/U1  ( .x(h[10]), .a(n5), .b(h[10]), .c(n3), .d(i[10]), 
        .e(\U10/nl ) );
    inv_1 \U9/Uii  ( .x(\U9/ni ), .a(i[9]) );
    inv_1 \U9/Uih  ( .x(\U9/nh ), .a(h[9]) );
    inv_1 \U9/Uil  ( .x(\U9/nl ), .a(l[9]) );
    ao23_1 \U9/Ucl/U1/U1  ( .x(l[9]), .a(n5), .b(l[9]), .c(n3), .d(\U9/ni ), 
        .e(\U9/nh ) );
    ao23_1 \U9/Uch/U1/U1  ( .x(h[9]), .a(n5), .b(h[9]), .c(n3), .d(i[9]), .e(
        \U9/nl ) );
    inv_1 \U8/Uii  ( .x(\U8/ni ), .a(i[8]) );
    inv_1 \U8/Uih  ( .x(\U8/nh ), .a(h[8]) );
    inv_1 \U8/Uil  ( .x(\U8/nl ), .a(l[8]) );
    ao23_1 \U8/Ucl/U1/U1  ( .x(l[8]), .a(n5), .b(l[8]), .c(n3), .d(\U8/ni ), 
        .e(\U8/nh ) );
    ao23_1 \U8/Uch/U1/U1  ( .x(h[8]), .a(n5), .b(h[8]), .c(n3), .d(i[8]), .e(
        \U8/nl ) );
    inv_1 \U7/Uii  ( .x(\U7/ni ), .a(i[7]) );
    inv_1 \U7/Uih  ( .x(\U7/nh ), .a(h[7]) );
    inv_1 \U7/Uil  ( .x(\U7/nl ), .a(l[7]) );
    ao23_1 \U7/Ucl/U1/U1  ( .x(l[7]), .a(n7), .b(l[7]), .c(n3), .d(\U7/ni ), 
        .e(\U7/nh ) );
    ao23_1 \U7/Uch/U1/U1  ( .x(h[7]), .a(n7), .b(h[7]), .c(n2), .d(i[7]), .e(
        \U7/nl ) );
    inv_1 \U6/Uii  ( .x(\U6/ni ), .a(i[6]) );
    inv_1 \U6/Uih  ( .x(\U6/nh ), .a(h[6]) );
    inv_1 \U6/Uil  ( .x(\U6/nl ), .a(l[6]) );
    ao23_1 \U6/Ucl/U1/U1  ( .x(l[6]), .a(n7), .b(l[6]), .c(n2), .d(\U6/ni ), 
        .e(\U6/nh ) );
    ao23_1 \U6/Uch/U1/U1  ( .x(h[6]), .a(n7), .b(h[6]), .c(n2), .d(i[6]), .e(
        \U6/nl ) );
    inv_1 \U5/Uii  ( .x(\U5/ni ), .a(i[5]) );
    inv_1 \U5/Uih  ( .x(\U5/nh ), .a(h[5]) );
    inv_1 \U5/Uil  ( .x(\U5/nl ), .a(l[5]) );
    ao23_1 \U5/Ucl/U1/U1  ( .x(l[5]), .a(n7), .b(l[5]), .c(n2), .d(\U5/ni ), 
        .e(\U5/nh ) );
    ao23_1 \U5/Uch/U1/U1  ( .x(h[5]), .a(n7), .b(h[5]), .c(n2), .d(i[5]), .e(
        \U5/nl ) );
    inv_1 \U4/Uii  ( .x(\U4/ni ), .a(i[4]) );
    inv_1 \U4/Uih  ( .x(\U4/nh ), .a(h[4]) );
    inv_1 \U4/Uil  ( .x(\U4/nl ), .a(l[4]) );
    ao23_1 \U4/Ucl/U1/U1  ( .x(l[4]), .a(n6), .b(l[4]), .c(n2), .d(\U4/ni ), 
        .e(\U4/nh ) );
    ao23_1 \U4/Uch/U1/U1  ( .x(h[4]), .a(n6), .b(h[4]), .c(n2), .d(i[4]), .e(
        \U4/nl ) );
    inv_1 \U3/Uii  ( .x(\U3/ni ), .a(i[3]) );
    inv_1 \U3/Uih  ( .x(\U3/nh ), .a(h[3]) );
    inv_1 \U3/Uil  ( .x(\U3/nl ), .a(l[3]) );
    ao23_1 \U3/Ucl/U1/U1  ( .x(l[3]), .a(n6), .b(l[3]), .c(n2), .d(\U3/ni ), 
        .e(\U3/nh ) );
    ao23_1 \U3/Uch/U1/U1  ( .x(h[3]), .a(n8), .b(h[3]), .c(n1), .d(i[3]), .e(
        \U3/nl ) );
    inv_1 \U2/Uii  ( .x(\U2/ni ), .a(i[2]) );
    inv_1 \U2/Uih  ( .x(\U2/nh ), .a(h[2]) );
    inv_1 \U2/Uil  ( .x(\U2/nl ), .a(l[2]) );
    ao23_1 \U2/Ucl/U1/U1  ( .x(l[2]), .a(n8), .b(l[2]), .c(n1), .d(\U2/ni ), 
        .e(\U2/nh ) );
    ao23_1 \U2/Uch/U1/U1  ( .x(h[2]), .a(n8), .b(h[2]), .c(n1), .d(i[2]), .e(
        \U2/nl ) );
    inv_1 \U1/Uii  ( .x(\U1/ni ), .a(i[1]) );
    inv_1 \U1/Uih  ( .x(\U1/nh ), .a(h[1]) );
    inv_1 \U1/Uil  ( .x(\U1/nl ), .a(l[1]) );
    ao23_1 \U1/Ucl/U1/U1  ( .x(l[1]), .a(n8), .b(l[1]), .c(n1), .d(\U1/ni ), 
        .e(\U1/nh ) );
    ao23_1 \U1/Uch/U1/U1  ( .x(h[1]), .a(n8), .b(h[1]), .c(n1), .d(i[1]), .e(
        \U1/nl ) );
    inv_1 \U0/Uii  ( .x(\U0/ni ), .a(i[0]) );
    inv_1 \U0/Uih  ( .x(\U0/nh ), .a(h[0]) );
    inv_1 \U0/Uil  ( .x(\U0/nl ), .a(l[0]) );
    ao23_1 \U0/Ucl/U1/U1  ( .x(l[0]), .a(n8), .b(l[0]), .c(n1), .d(\U0/ni ), 
        .e(\U0/nh ) );
    ao23_1 \U0/Uch/U1/U1  ( .x(h[0]), .a(n8), .b(h[0]), .c(n1), .d(i[0]), .e(
        \U0/nl ) );
    buf_16 U1 ( .x(n1), .a(n12) );
    buf_16 U2 ( .x(n2), .a(n12) );
    buf_16 U3 ( .x(n3), .a(n12) );
    buf_16 U4 ( .x(n4), .a(n11) );
    buf_16 U5 ( .x(n5), .a(n11) );
    buf_16 U6 ( .x(n6), .a(n11) );
    buf_16 U7 ( .x(n7), .a(n10) );
    buf_16 U8 ( .x(n8), .a(n10) );
    buf_16 U9 ( .x(n9), .a(n10) );
    buf_16 U10 ( .x(n10), .a(req) );
    buf_16 U11 ( .x(n11), .a(req) );
    buf_16 U12 ( .x(n12), .a(req) );
endmodule


module sr2dr_word_3 ( i, req, h, l );
input  [31:0] i;
output [31:0] h;
output [31:0] l;
input  req;
    wire \U31/nl , \U31/ni , \U31/nh , \U30/nl , \U30/ni , \U30/nh , \U29/nl , 
        \U29/ni , \U29/nh , \U28/nl , \U28/ni , \U28/nh , \U27/nl , \U27/ni , 
        \U27/nh , \U26/nl , \U26/ni , \U26/nh , \U25/nl , \U25/ni , \U25/nh , 
        \U24/nl , \U24/ni , \U24/nh , \U23/nl , \U23/ni , \U23/nh , \U22/nl , 
        \U22/ni , \U22/nh , \U21/nl , \U21/ni , \U21/nh , \U20/nl , \U20/ni , 
        \U20/nh , \U19/nl , \U19/ni , \U19/nh , \U18/nl , \U18/ni , \U18/nh , 
        \U17/nl , \U17/ni , \U17/nh , \U16/nl , \U16/ni , \U16/nh , \U15/nl , 
        \U15/ni , \U15/nh , \U14/nl , \U14/ni , \U14/nh , \U13/nl , \U13/ni , 
        \U13/nh , \U12/nl , \U12/ni , \U12/nh , \U11/nl , \U11/ni , \U11/nh , 
        \U10/nl , \U10/ni , \U10/nh , \U9/nl , \U9/ni , \U9/nh , \U8/nl , 
        \U8/ni , \U8/nh , \U7/nl , \U7/ni , \U7/nh , \U6/nl , \U6/ni , \U6/nh , 
        \U5/nl , \U5/ni , \U5/nh , \U4/nl , \U4/ni , \U4/nh , \U3/nl , \U3/ni , 
        \U3/nh , \U2/nl , \U2/ni , \U2/nh , \U1/nl , \U1/ni , \U1/nh , \U0/nl , 
        \U0/ni , \U0/nh , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
    inv_1 \U31/Uii  ( .x(\U31/ni ), .a(i[31]) );
    inv_1 \U31/Uih  ( .x(\U31/nh ), .a(h[31]) );
    inv_1 \U31/Uil  ( .x(\U31/nl ), .a(l[31]) );
    ao23_1 \U31/Ucl/U1/U1  ( .x(l[31]), .a(n9), .b(l[31]), .c(n1), .d(\U31/ni 
        ), .e(\U31/nh ) );
    ao23_1 \U31/Uch/U1/U1  ( .x(h[31]), .a(n9), .b(h[31]), .c(n2), .d(i[31]), 
        .e(\U31/nl ) );
    inv_1 \U30/Uii  ( .x(\U30/ni ), .a(i[30]) );
    inv_1 \U30/Uih  ( .x(\U30/nh ), .a(h[30]) );
    inv_1 \U30/Uil  ( .x(\U30/nl ), .a(l[30]) );
    ao23_1 \U30/Ucl/U1/U1  ( .x(l[30]), .a(n8), .b(l[30]), .c(n1), .d(\U30/ni 
        ), .e(\U30/nh ) );
    ao23_1 \U30/Uch/U1/U1  ( .x(h[30]), .a(n8), .b(h[30]), .c(n1), .d(i[30]), 
        .e(\U30/nl ) );
    inv_1 \U29/Uii  ( .x(\U29/ni ), .a(i[29]) );
    inv_1 \U29/Uih  ( .x(\U29/nh ), .a(h[29]) );
    inv_1 \U29/Uil  ( .x(\U29/nl ), .a(l[29]) );
    ao23_1 \U29/Ucl/U1/U1  ( .x(l[29]), .a(n8), .b(l[29]), .c(n1), .d(\U29/ni 
        ), .e(\U29/nh ) );
    ao23_1 \U29/Uch/U1/U1  ( .x(h[29]), .a(n8), .b(h[29]), .c(n2), .d(i[29]), 
        .e(\U29/nl ) );
    inv_1 \U28/Uii  ( .x(\U28/ni ), .a(i[28]) );
    inv_1 \U28/Uih  ( .x(\U28/nh ), .a(h[28]) );
    inv_1 \U28/Uil  ( .x(\U28/nl ), .a(l[28]) );
    ao23_1 \U28/Ucl/U1/U1  ( .x(l[28]), .a(n8), .b(l[28]), .c(n2), .d(\U28/ni 
        ), .e(\U28/nh ) );
    ao23_1 \U28/Uch/U1/U1  ( .x(h[28]), .a(n8), .b(h[28]), .c(n2), .d(i[28]), 
        .e(\U28/nl ) );
    inv_1 \U27/Uii  ( .x(\U27/ni ), .a(i[27]) );
    inv_1 \U27/Uih  ( .x(\U27/nh ), .a(h[27]) );
    inv_1 \U27/Uil  ( .x(\U27/nl ), .a(l[27]) );
    ao23_1 \U27/Ucl/U1/U1  ( .x(l[27]), .a(n8), .b(l[27]), .c(n2), .d(\U27/ni 
        ), .e(\U27/nh ) );
    ao23_1 \U27/Uch/U1/U1  ( .x(h[27]), .a(n8), .b(h[27]), .c(n2), .d(i[27]), 
        .e(\U27/nl ) );
    inv_1 \U26/Uii  ( .x(\U26/ni ), .a(i[26]) );
    inv_1 \U26/Uih  ( .x(\U26/nh ), .a(h[26]) );
    inv_1 \U26/Uil  ( .x(\U26/nl ), .a(l[26]) );
    ao23_1 \U26/Ucl/U1/U1  ( .x(l[26]), .a(n7), .b(l[26]), .c(n2), .d(\U26/ni 
        ), .e(\U26/nh ) );
    ao23_1 \U26/Uch/U1/U1  ( .x(h[26]), .a(n7), .b(h[26]), .c(n4), .d(i[26]), 
        .e(\U26/nl ) );
    inv_1 \U25/Uii  ( .x(\U25/ni ), .a(i[25]) );
    inv_1 \U25/Uih  ( .x(\U25/nh ), .a(h[25]) );
    inv_1 \U25/Uil  ( .x(\U25/nl ), .a(l[25]) );
    ao23_1 \U25/Ucl/U1/U1  ( .x(l[25]), .a(n7), .b(l[25]), .c(n4), .d(\U25/ni 
        ), .e(\U25/nh ) );
    ao23_1 \U25/Uch/U1/U1  ( .x(h[25]), .a(n7), .b(h[25]), .c(n4), .d(i[25]), 
        .e(\U25/nl ) );
    inv_1 \U24/Uii  ( .x(\U24/ni ), .a(i[24]) );
    inv_1 \U24/Uih  ( .x(\U24/nh ), .a(h[24]) );
    inv_1 \U24/Uil  ( .x(\U24/nl ), .a(l[24]) );
    ao23_1 \U24/Ucl/U1/U1  ( .x(l[24]), .a(n7), .b(l[24]), .c(n4), .d(\U24/ni 
        ), .e(\U24/nh ) );
    ao23_1 \U24/Uch/U1/U1  ( .x(h[24]), .a(n7), .b(h[24]), .c(n4), .d(i[24]), 
        .e(\U24/nl ) );
    inv_1 \U23/Uii  ( .x(\U23/ni ), .a(i[23]) );
    inv_1 \U23/Uih  ( .x(\U23/nh ), .a(h[23]) );
    inv_1 \U23/Uil  ( .x(\U23/nl ), .a(l[23]) );
    ao23_1 \U23/Ucl/U1/U1  ( .x(l[23]), .a(n7), .b(l[23]), .c(n3), .d(\U23/ni 
        ), .e(\U23/nh ) );
    ao23_1 \U23/Uch/U1/U1  ( .x(h[23]), .a(n7), .b(h[23]), .c(n3), .d(i[23]), 
        .e(\U23/nl ) );
    inv_1 \U22/Uii  ( .x(\U22/ni ), .a(i[22]) );
    inv_1 \U22/Uih  ( .x(\U22/nh ), .a(h[22]) );
    inv_1 \U22/Uil  ( .x(\U22/nl ), .a(l[22]) );
    ao23_1 \U22/Ucl/U1/U1  ( .x(l[22]), .a(n6), .b(l[22]), .c(n3), .d(\U22/ni 
        ), .e(\U22/nh ) );
    ao23_1 \U22/Uch/U1/U1  ( .x(h[22]), .a(n6), .b(h[22]), .c(n3), .d(i[22]), 
        .e(\U22/nl ) );
    inv_1 \U21/Uii  ( .x(\U21/ni ), .a(i[21]) );
    inv_1 \U21/Uih  ( .x(\U21/nh ), .a(h[21]) );
    inv_1 \U21/Uil  ( .x(\U21/nl ), .a(l[21]) );
    ao23_1 \U21/Ucl/U1/U1  ( .x(l[21]), .a(n6), .b(l[21]), .c(n3), .d(\U21/ni 
        ), .e(\U21/nh ) );
    ao23_1 \U21/Uch/U1/U1  ( .x(h[21]), .a(n6), .b(h[21]), .c(n3), .d(i[21]), 
        .e(\U21/nl ) );
    inv_1 \U20/Uii  ( .x(\U20/ni ), .a(i[20]) );
    inv_1 \U20/Uih  ( .x(\U20/nh ), .a(h[20]) );
    inv_1 \U20/Uil  ( .x(\U20/nl ), .a(l[20]) );
    ao23_1 \U20/Ucl/U1/U1  ( .x(l[20]), .a(n6), .b(l[20]), .c(n5), .d(\U20/ni 
        ), .e(\U20/nh ) );
    ao23_1 \U20/Uch/U1/U1  ( .x(h[20]), .a(n6), .b(h[20]), .c(n4), .d(i[20]), 
        .e(\U20/nl ) );
    inv_1 \U19/Uii  ( .x(\U19/ni ), .a(i[19]) );
    inv_1 \U19/Uih  ( .x(\U19/nh ), .a(h[19]) );
    inv_1 \U19/Uil  ( .x(\U19/nl ), .a(l[19]) );
    ao23_1 \U19/Ucl/U1/U1  ( .x(l[19]), .a(n6), .b(l[19]), .c(n4), .d(\U19/ni 
        ), .e(\U19/nh ) );
    ao23_1 \U19/Uch/U1/U1  ( .x(h[19]), .a(n6), .b(h[19]), .c(n4), .d(i[19]), 
        .e(\U19/nl ) );
    inv_1 \U18/Uii  ( .x(\U18/ni ), .a(i[18]) );
    inv_1 \U18/Uih  ( .x(\U18/nh ), .a(h[18]) );
    inv_1 \U18/Uil  ( .x(\U18/nl ), .a(l[18]) );
    ao23_1 \U18/Ucl/U1/U1  ( .x(l[18]), .a(n5), .b(l[18]), .c(n5), .d(\U18/ni 
        ), .e(\U18/nh ) );
    ao23_1 \U18/Uch/U1/U1  ( .x(h[18]), .a(n5), .b(h[18]), .c(n5), .d(i[18]), 
        .e(\U18/nl ) );
    inv_1 \U17/Uii  ( .x(\U17/ni ), .a(i[17]) );
    inv_1 \U17/Uih  ( .x(\U17/nh ), .a(h[17]) );
    inv_1 \U17/Uil  ( .x(\U17/nl ), .a(l[17]) );
    ao23_1 \U17/Ucl/U1/U1  ( .x(l[17]), .a(n6), .b(l[17]), .c(n5), .d(\U17/ni 
        ), .e(\U17/nh ) );
    ao23_1 \U17/Uch/U1/U1  ( .x(h[17]), .a(n7), .b(h[17]), .c(n4), .d(i[17]), 
        .e(\U17/nl ) );
    inv_1 \U16/Uii  ( .x(\U16/ni ), .a(i[16]) );
    inv_1 \U16/Uih  ( .x(\U16/nh ), .a(h[16]) );
    inv_1 \U16/Uil  ( .x(\U16/nl ), .a(l[16]) );
    ao23_1 \U16/Ucl/U1/U1  ( .x(l[16]), .a(n9), .b(l[16]), .c(n3), .d(\U16/ni 
        ), .e(\U16/nh ) );
    ao23_1 \U16/Uch/U1/U1  ( .x(h[16]), .a(n9), .b(h[16]), .c(n1), .d(i[16]), 
        .e(\U16/nl ) );
    inv_1 \U15/Uii  ( .x(\U15/ni ), .a(i[15]) );
    inv_1 \U15/Uih  ( .x(\U15/nh ), .a(h[15]) );
    inv_1 \U15/Uil  ( .x(\U15/nl ), .a(l[15]) );
    ao23_1 \U15/Ucl/U1/U1  ( .x(l[15]), .a(n8), .b(l[15]), .c(n1), .d(\U15/ni 
        ), .e(\U15/nh ) );
    ao23_1 \U15/Uch/U1/U1  ( .x(h[15]), .a(n7), .b(h[15]), .c(n1), .d(i[15]), 
        .e(\U15/nl ) );
    inv_1 \U14/Uii  ( .x(\U14/ni ), .a(i[14]) );
    inv_1 \U14/Uih  ( .x(\U14/nh ), .a(h[14]) );
    inv_1 \U14/Uil  ( .x(\U14/nl ), .a(l[14]) );
    ao23_1 \U14/Ucl/U1/U1  ( .x(l[14]), .a(n6), .b(l[14]), .c(n1), .d(\U14/ni 
        ), .e(\U14/nh ) );
    ao23_1 \U14/Uch/U1/U1  ( .x(h[14]), .a(n6), .b(h[14]), .c(n3), .d(i[14]), 
        .e(\U14/nl ) );
    inv_1 \U13/Uii  ( .x(\U13/ni ), .a(i[13]) );
    inv_1 \U13/Uih  ( .x(\U13/nh ), .a(h[13]) );
    inv_1 \U13/Uil  ( .x(\U13/nl ), .a(l[13]) );
    ao23_1 \U13/Ucl/U1/U1  ( .x(l[13]), .a(n6), .b(l[13]), .c(n4), .d(\U13/ni 
        ), .e(\U13/nh ) );
    ao23_1 \U13/Uch/U1/U1  ( .x(h[13]), .a(n6), .b(h[13]), .c(n4), .d(i[13]), 
        .e(\U13/nl ) );
    inv_1 \U12/Uii  ( .x(\U12/ni ), .a(i[12]) );
    inv_1 \U12/Uih  ( .x(\U12/nh ), .a(h[12]) );
    inv_1 \U12/Uil  ( .x(\U12/nl ), .a(l[12]) );
    ao23_1 \U12/Ucl/U1/U1  ( .x(l[12]), .a(n5), .b(l[12]), .c(n4), .d(\U12/ni 
        ), .e(\U12/nh ) );
    ao23_1 \U12/Uch/U1/U1  ( .x(h[12]), .a(n5), .b(h[12]), .c(n4), .d(i[12]), 
        .e(\U12/nl ) );
    inv_1 \U11/Uii  ( .x(\U11/ni ), .a(i[11]) );
    inv_1 \U11/Uih  ( .x(\U11/nh ), .a(h[11]) );
    inv_1 \U11/Uil  ( .x(\U11/nl ), .a(l[11]) );
    ao23_1 \U11/Ucl/U1/U1  ( .x(l[11]), .a(n5), .b(l[11]), .c(n4), .d(\U11/ni 
        ), .e(\U11/nh ) );
    ao23_1 \U11/Uch/U1/U1  ( .x(h[11]), .a(n5), .b(h[11]), .c(n4), .d(i[11]), 
        .e(\U11/nl ) );
    inv_1 \U10/Uii  ( .x(\U10/ni ), .a(i[10]) );
    inv_1 \U10/Uih  ( .x(\U10/nh ), .a(h[10]) );
    inv_1 \U10/Uil  ( .x(\U10/nl ), .a(l[10]) );
    ao23_1 \U10/Ucl/U1/U1  ( .x(l[10]), .a(n5), .b(l[10]), .c(n3), .d(\U10/ni 
        ), .e(\U10/nh ) );
    ao23_1 \U10/Uch/U1/U1  ( .x(h[10]), .a(n5), .b(h[10]), .c(n3), .d(i[10]), 
        .e(\U10/nl ) );
    inv_1 \U9/Uii  ( .x(\U9/ni ), .a(i[9]) );
    inv_1 \U9/Uih  ( .x(\U9/nh ), .a(h[9]) );
    inv_1 \U9/Uil  ( .x(\U9/nl ), .a(l[9]) );
    ao23_1 \U9/Ucl/U1/U1  ( .x(l[9]), .a(n5), .b(l[9]), .c(n3), .d(\U9/ni ), 
        .e(\U9/nh ) );
    ao23_1 \U9/Uch/U1/U1  ( .x(h[9]), .a(n5), .b(h[9]), .c(n3), .d(i[9]), .e(
        \U9/nl ) );
    inv_1 \U8/Uii  ( .x(\U8/ni ), .a(i[8]) );
    inv_1 \U8/Uih  ( .x(\U8/nh ), .a(h[8]) );
    inv_1 \U8/Uil  ( .x(\U8/nl ), .a(l[8]) );
    ao23_1 \U8/Ucl/U1/U1  ( .x(l[8]), .a(n5), .b(l[8]), .c(n3), .d(\U8/ni ), 
        .e(\U8/nh ) );
    ao23_1 \U8/Uch/U1/U1  ( .x(h[8]), .a(n5), .b(h[8]), .c(n3), .d(i[8]), .e(
        \U8/nl ) );
    inv_1 \U7/Uii  ( .x(\U7/ni ), .a(i[7]) );
    inv_1 \U7/Uih  ( .x(\U7/nh ), .a(h[7]) );
    inv_1 \U7/Uil  ( .x(\U7/nl ), .a(l[7]) );
    ao23_1 \U7/Ucl/U1/U1  ( .x(l[7]), .a(n7), .b(l[7]), .c(n3), .d(\U7/ni ), 
        .e(\U7/nh ) );
    ao23_1 \U7/Uch/U1/U1  ( .x(h[7]), .a(n7), .b(h[7]), .c(n2), .d(i[7]), .e(
        \U7/nl ) );
    inv_1 \U6/Uii  ( .x(\U6/ni ), .a(i[6]) );
    inv_1 \U6/Uih  ( .x(\U6/nh ), .a(h[6]) );
    inv_1 \U6/Uil  ( .x(\U6/nl ), .a(l[6]) );
    ao23_1 \U6/Ucl/U1/U1  ( .x(l[6]), .a(n7), .b(l[6]), .c(n2), .d(\U6/ni ), 
        .e(\U6/nh ) );
    ao23_1 \U6/Uch/U1/U1  ( .x(h[6]), .a(n7), .b(h[6]), .c(n2), .d(i[6]), .e(
        \U6/nl ) );
    inv_1 \U5/Uii  ( .x(\U5/ni ), .a(i[5]) );
    inv_1 \U5/Uih  ( .x(\U5/nh ), .a(h[5]) );
    inv_1 \U5/Uil  ( .x(\U5/nl ), .a(l[5]) );
    ao23_1 \U5/Ucl/U1/U1  ( .x(l[5]), .a(n7), .b(l[5]), .c(n2), .d(\U5/ni ), 
        .e(\U5/nh ) );
    ao23_1 \U5/Uch/U1/U1  ( .x(h[5]), .a(n7), .b(h[5]), .c(n2), .d(i[5]), .e(
        \U5/nl ) );
    inv_1 \U4/Uii  ( .x(\U4/ni ), .a(i[4]) );
    inv_1 \U4/Uih  ( .x(\U4/nh ), .a(h[4]) );
    inv_1 \U4/Uil  ( .x(\U4/nl ), .a(l[4]) );
    ao23_1 \U4/Ucl/U1/U1  ( .x(l[4]), .a(n6), .b(l[4]), .c(n2), .d(\U4/ni ), 
        .e(\U4/nh ) );
    ao23_1 \U4/Uch/U1/U1  ( .x(h[4]), .a(n6), .b(h[4]), .c(n2), .d(i[4]), .e(
        \U4/nl ) );
    inv_1 \U3/Uii  ( .x(\U3/ni ), .a(i[3]) );
    inv_1 \U3/Uih  ( .x(\U3/nh ), .a(h[3]) );
    inv_1 \U3/Uil  ( .x(\U3/nl ), .a(l[3]) );
    ao23_1 \U3/Ucl/U1/U1  ( .x(l[3]), .a(n6), .b(l[3]), .c(n2), .d(\U3/ni ), 
        .e(\U3/nh ) );
    ao23_1 \U3/Uch/U1/U1  ( .x(h[3]), .a(n8), .b(h[3]), .c(n1), .d(i[3]), .e(
        \U3/nl ) );
    inv_1 \U2/Uii  ( .x(\U2/ni ), .a(i[2]) );
    inv_1 \U2/Uih  ( .x(\U2/nh ), .a(h[2]) );
    inv_1 \U2/Uil  ( .x(\U2/nl ), .a(l[2]) );
    ao23_1 \U2/Ucl/U1/U1  ( .x(l[2]), .a(n8), .b(l[2]), .c(n1), .d(\U2/ni ), 
        .e(\U2/nh ) );
    ao23_1 \U2/Uch/U1/U1  ( .x(h[2]), .a(n8), .b(h[2]), .c(n1), .d(i[2]), .e(
        \U2/nl ) );
    inv_1 \U1/Uii  ( .x(\U1/ni ), .a(i[1]) );
    inv_1 \U1/Uih  ( .x(\U1/nh ), .a(h[1]) );
    inv_1 \U1/Uil  ( .x(\U1/nl ), .a(l[1]) );
    ao23_1 \U1/Ucl/U1/U1  ( .x(l[1]), .a(n8), .b(l[1]), .c(n1), .d(\U1/ni ), 
        .e(\U1/nh ) );
    ao23_1 \U1/Uch/U1/U1  ( .x(h[1]), .a(n8), .b(h[1]), .c(n1), .d(i[1]), .e(
        \U1/nl ) );
    inv_1 \U0/Uii  ( .x(\U0/ni ), .a(i[0]) );
    inv_1 \U0/Uih  ( .x(\U0/nh ), .a(h[0]) );
    inv_1 \U0/Uil  ( .x(\U0/nl ), .a(l[0]) );
    ao23_1 \U0/Ucl/U1/U1  ( .x(l[0]), .a(n8), .b(l[0]), .c(n1), .d(\U0/ni ), 
        .e(\U0/nh ) );
    ao23_1 \U0/Uch/U1/U1  ( .x(h[0]), .a(n8), .b(h[0]), .c(n1), .d(i[0]), .e(
        \U0/nl ) );
    buf_16 U1 ( .x(n1), .a(n12) );
    buf_16 U2 ( .x(n2), .a(n12) );
    buf_16 U3 ( .x(n3), .a(n12) );
    buf_16 U4 ( .x(n4), .a(n11) );
    buf_16 U5 ( .x(n5), .a(n11) );
    buf_16 U6 ( .x(n6), .a(n11) );
    buf_16 U7 ( .x(n7), .a(n10) );
    buf_16 U8 ( .x(n8), .a(n10) );
    buf_16 U9 ( .x(n9), .a(n10) );
    buf_16 U10 ( .x(n10), .a(req) );
    buf_16 U11 ( .x(n11), .a(req) );
    buf_16 U12 ( .x(n12), .a(req) );
endmodule


module latch_ctrl_1 ( rin, ain, rout, aout, en, reset );
input  rin, aout, reset;
output ain, rout, en;
    wire N5, N6, na, a, n_rout, nreset, n3, \c_rout/ob , n1;
    inv_1 U0 ( .x(nreset), .a(reset) );
    nor2_1 U1 ( .x(ain), .a(na), .b(n1) );
    inv_1 U2 ( .x(na), .a(a) );
    inv_1 U3 ( .x(N6), .a(N5) );
    inv_1 U4 ( .x(rout), .a(n_rout) );
    and2_1 C9 ( .x(n3), .a(na), .b(N6) );
    or2_1 C11 ( .x(N5), .a(rout), .b(aout) );
    oa21_1 \c_na/__tmp99/U1  ( .x(a), .a(n1), .b(a), .c(rin) );
    oai21_1 \c_rout/U1  ( .x(\c_rout/ob ), .a(aout), .b(n_rout), .c(na) );
    nand2_1 \c_rout/U2  ( .x(n_rout), .a(nreset), .b(\c_rout/ob ) );
    buf_1 U5 ( .x(en), .a(n3) );
    buf_1 U6 ( .x(n1), .a(n3) );
endmodule


module m2cp_dport ( req_in, ts_o, sel_o, mult_o, we_o, prd_o, seq_o, adr_o, 
    dat_o, ain, ic_seq, ic_pred, ic_size, ic_itag, ic_wd, ic_lock, ic_a, 
    ic_rnw, ic_col, ic_ack, req_out, ts_i, we_i, err_i, rty_i, acc_i, dat_i, 
    aout, ir_rd, ir_err, ir_rnw, ir_ack, tag_id, reset );
input  [2:0] ts_o;
input  [3:0] sel_o;
input  [31:0] adr_o;
input  [31:0] dat_o;
output [1:0] ic_seq;
output [1:0] ic_pred;
output [3:0] ic_size;
output [9:0] ic_itag;
output [63:0] ic_wd;
output [1:0] ic_lock;
output [63:0] ic_a;
output [1:0] ic_rnw;
output [5:0] ic_col;
output [2:0] ts_i;
output [31:0] dat_i;
input  [63:0] ir_rd;
input  [1:0] ir_err;
input  [1:0] ir_rnw;
input  [4:0] tag_id;
input  req_in, mult_o, we_o, prd_o, seq_o, ic_ack, aout, reset;
output ain, req_out, we_i, err_i, rty_i, acc_i, ir_ack;
    wire n63, n64, n65, n68, n69, n70, n72, n73, n74, n75, n76, n77, n78, n79, 
        n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, 
        n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, 
        n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
        n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, 
        n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
        n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
        n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
        n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
        n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
        n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, 
        n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, 
        n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, 
        n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, 
        n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, 
        n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, 
        n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, 
        n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, 
        n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, 
        n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n2, n3, n4, 
        n5, req_in_delayed, \size[1] , \size[0] , \data[15] , \data[14] , 
        \data[13] , \data[12] , \data[11] , \data[10] , \data[9] , \data[8] , 
        \data[7] , \data[6] , \data[5] , \data[4] , \data[3] , \data[2] , 
        \data[1] , \data[0] , _24_net_, _25_net_, _26_net_, comp_basic, 
        high_ir_rd, low_ir_rd, comp_rd, _27_net_, all_r, _28_net_, all_w, 
        complete, complete_delayed, en, \all_read/__tmp99/loop , \Ucol2/nl , 
        \Ucol2/ni , \Ucol2/nh , \Ucol1/nl , \Ucol1/ni , \Ucol1/nh , \Ucol0/nl , 
        \Ucol0/ni , \Ucol0/nh , \Utag4/nl , \Utag4/ni , \Utag4/nh , \Utag3/nl , 
        \Utag3/ni , \Utag3/nh , \Utag2/nl , \Utag2/ni , \Utag2/nh , \Utag1/nl , 
        \Utag1/ni , \Utag1/nh , \Utag0/nl , \Utag0/ni , \Utag0/nh , \Usze1/nl , 
        \Usze1/ni , \Usze1/nh , \Usze0/nl , \Usze0/ni , \Usze0/nh , \Urnw/nl , 
        \Urnw/ni , \Urnw/nh , \Ulock/nl , \Ulock/ni , \Ulock/nh , \Upred/nl , 
        \Upred/ni , \Upred/nh , \Useq/nl , \Useq/ni , \Useq/nh , n1, n6, n7, 
        n8, n9, n10, n11;
    assign ain = ic_ack;
    assign ts_i[2] = 1'b0;
    assign ts_i[1] = 1'b0;
    assign ts_i[0] = 1'b0;
    assign rty_i = 1'b0;
    assign acc_i = 1'b0;
    matched_delay_m2cp_com_dport U130 ( .x(req_in_delayed), .a(req_in) );
    sr2dr_word_3 Uwd ( .i({dat_o[31], dat_o[30], dat_o[29], dat_o[28], 
        dat_o[27], dat_o[26], dat_o[25], dat_o[24], dat_o[23], dat_o[22], 
        dat_o[21], dat_o[20], dat_o[19], dat_o[18], dat_o[17], dat_o[16], 
        \data[15] , \data[14] , \data[13] , \data[12] , \data[11] , \data[10] , 
        \data[9] , \data[8] , \data[7] , \data[6] , \data[5] , \data[4] , 
        \data[3] , \data[2] , \data[1] , \data[0] }), .req(n8), .h(ic_wd
        [63:32]), .l(ic_wd[31:0]) );
    sr2dr_word_2 Ua ( .i(adr_o), .req(n8), .h(ic_a[63:32]), .l(ic_a[31:0]) );
    latch_ctrl_1 lc ( .rin(complete_delayed), .ain(ir_ack), .rout(req_out), 
        .aout(aout), .en(en), .reset(reset) );
    nand2i_1 U59 ( .x(_28_net_), .a(ir_err[1]), .b(n72) );
    nand2_1 U61 ( .x(_26_net_), .a(n72), .b(n77) );
    nand2i_1 U112 ( .x(_25_net_), .a(ir_err[1]), .b(n78) );
    and2_1 U274 ( .x(_27_net_), .a(ir_rnw[1]), .b(ir_err[0]) );
    inv_1 U275 ( .x(_24_net_), .a(we_o) );
    inv_1 U2 ( .x(n112), .a(ir_rd[4]) );
    inv_1 U3 ( .x(n124), .a(ir_rd[0]) );
    inv_1 U4 ( .x(n118), .a(ir_rd[2]) );
    inv_1 U5 ( .x(n206), .a(dat_o[28]) );
    inv_1 U6 ( .x(n208), .a(dat_o[27]) );
    inv_1 U7 ( .x(n210), .a(dat_o[26]) );
    inv_1 U8 ( .x(n197), .a(dat_o[25]) );
    inv_1 U9 ( .x(n199), .a(dat_o[24]) );
    inv_1 U10 ( .x(n202), .a(dat_o[15]) );
    inv_1 U11 ( .x(n201), .a(dat_o[31]) );
    inv_1 U12 ( .x(n203), .a(dat_o[30]) );
    inv_1 U13 ( .x(n204), .a(dat_o[29]) );
    nor2_1 U14 ( .x(\size[1] ), .a(n83), .b(n84) );
    inv_1 U15 ( .x(n72), .a(ir_rnw[0]) );
    oa21_1 U16 ( .x(n89), .a(n205), .b(n64), .c(n2) );
    inv_1 U24 ( .x(n2), .a(n90) );
    inv_1 U17 ( .x(n205), .a(dat_o[13]) );
    inv_1 U18 ( .x(n64), .a(sel_o[1]) );
    oa21_1 U19 ( .x(n97), .a(n198), .b(n64), .c(n3) );
    inv_1 U276 ( .x(n3), .a(n98) );
    inv_1 U20 ( .x(n198), .a(dat_o[9]) );
    oa21_1 U21 ( .x(n87), .a(n63), .b(n64), .c(n4) );
    inv_1 U277 ( .x(n4), .a(n88) );
    inv_1 U22 ( .x(n63), .a(dat_o[14]) );
    oa21_1 U23 ( .x(n85), .a(n202), .b(n64), .c(n5) );
    inv_1 U278 ( .x(n5), .a(n86) );
    nand2_1 U25 ( .x(n290), .a(n289), .b(n288) );
    nand2_1 U26 ( .x(n79), .a(n277), .b(n270) );
    nor2_1 U27 ( .x(n277), .a(n273), .b(n276) );
    nor2_1 U28 ( .x(n270), .a(n266), .b(n269) );
    nand2_1 U29 ( .x(n283), .a(n282), .b(n281) );
    nand2_1 U30 ( .x(n298), .a(dat_o[20]), .b(n70) );
    inv_1 U31 ( .x(n70), .a(n68) );
    nand2_1 U32 ( .x(n213), .a(n223), .b(sel_o[1]) );
    nand2_1 U33 ( .x(n80), .a(n291), .b(n284) );
    nor2_1 U34 ( .x(n291), .a(n287), .b(n290) );
    nor2_1 U35 ( .x(n284), .a(n280), .b(n283) );
    aoi21_1 U36 ( .x(n99), .a(dat_o[8]), .b(sel_o[1]), .c(n100) );
    aoi21_1 U37 ( .x(n95), .a(dat_o[10]), .b(sel_o[1]), .c(n96) );
    aoi21_1 U38 ( .x(n93), .a(dat_o[11]), .b(sel_o[1]), .c(n94) );
    aoi21_1 U39 ( .x(n91), .a(dat_o[12]), .b(sel_o[1]), .c(n92) );
    inv_1 U40 ( .x(n81), .a(all_r) );
    nand2_1 U42 ( .x(n84), .a(sel_o[0]), .b(sel_o[1]) );
    inv_1 U45 ( .x(n68), .a(sel_o[2]) );
    inv_1 U46 ( .x(n69), .a(n68) );
    nand2_1 U48 ( .x(n83), .a(n70), .b(sel_o[3]) );
    nand2_1 U51 ( .x(n300), .a(dat_o[19]), .b(n69) );
    nand2_1 U52 ( .x(n294), .a(dat_o[22]), .b(n69) );
    nand2_1 U53 ( .x(n302), .a(dat_o[18]), .b(n69) );
    nand2_1 U54 ( .x(n296), .a(dat_o[21]), .b(n69) );
    nand2_1 U55 ( .x(n306), .a(dat_o[16]), .b(n69) );
    nand2_1 U56 ( .x(n292), .a(dat_o[23]), .b(n69) );
    nand2_1 U57 ( .x(n304), .a(dat_o[17]), .b(n69) );
    nand4_1 U60 ( .x(low_ir_rd), .a(n73), .b(n74), .c(n75), .d(n76) );
    nand2_1 U62 ( .x(complete), .a(n81), .b(n82) );
    matched_delay_m2cp_resp_dport mdel ( .x(complete_delayed), .a(complete) );
    inv_1 U63 ( .x(n200), .a(dat_o[8]) );
    inv_1 U64 ( .x(n207), .a(dat_o[12]) );
    inv_1 U65 ( .x(n209), .a(dat_o[11]) );
    inv_1 U66 ( .x(n211), .a(dat_o[10]) );
    nand4_1 U67 ( .x(n224), .a(n225), .b(n226), .c(n227), .d(n228) );
    nand4_1 U68 ( .x(n229), .a(n230), .b(n231), .c(n232), .d(n233) );
    nor2_1 U69 ( .x(n76), .a(n224), .b(n229) );
    nand4_1 U70 ( .x(n234), .a(n235), .b(n236), .c(n237), .d(n238) );
    nand4_1 U71 ( .x(n239), .a(n240), .b(n241), .c(n242), .d(n243) );
    nor2_1 U72 ( .x(n75), .a(n234), .b(n239) );
    nand4_1 U73 ( .x(n244), .a(n245), .b(n246), .c(n247), .d(n248) );
    nand4_1 U74 ( .x(n249), .a(n250), .b(n251), .c(n252), .d(n253) );
    nor2_1 U75 ( .x(n74), .a(n244), .b(n249) );
    nand4_1 U76 ( .x(n254), .a(n255), .b(n256), .c(n257), .d(n258) );
    nand4_1 U77 ( .x(n259), .a(n260), .b(n261), .c(n262), .d(n263) );
    nor2_1 U78 ( .x(n73), .a(n254), .b(n259) );
    nand2_1 U79 ( .x(n266), .a(n265), .b(n264) );
    nand2_1 U80 ( .x(n269), .a(n268), .b(n267) );
    nand2_1 U81 ( .x(n273), .a(n272), .b(n271) );
    nand2_1 U82 ( .x(n276), .a(n275), .b(n274) );
    nand2_1 U83 ( .x(n280), .a(n279), .b(n278) );
    nand2_1 U84 ( .x(n287), .a(n286), .b(n285) );
    nand2_1 U85 ( .x(n86), .a(n292), .b(n293) );
    nand2_1 U86 ( .x(n88), .a(n294), .b(n295) );
    nand2_1 U87 ( .x(n90), .a(n296), .b(n297) );
    nand2_1 U88 ( .x(n92), .a(n298), .b(n299) );
    nand2_1 U89 ( .x(n94), .a(n300), .b(n301) );
    nand2_1 U90 ( .x(n96), .a(n302), .b(n303) );
    nand2_1 U91 ( .x(n98), .a(n304), .b(n305) );
    nand2_1 U92 ( .x(n100), .a(n306), .b(n307) );
    inv_1 U93 ( .x(n222), .a(dat_o[0]) );
    inv_1 U94 ( .x(n221), .a(dat_o[1]) );
    inv_1 U95 ( .x(n220), .a(dat_o[2]) );
    inv_1 U96 ( .x(n219), .a(dat_o[3]) );
    inv_1 U97 ( .x(n218), .a(dat_o[4]) );
    inv_1 U98 ( .x(n217), .a(dat_o[5]) );
    inv_1 U99 ( .x(n216), .a(dat_o[6]) );
    inv_1 U100 ( .x(n215), .a(dat_o[7]) );
    inv_1 U101 ( .x(n77), .a(ir_rnw[1]) );
    inv_1 U103 ( .x(n82), .a(all_w) );
    nand2_1 U104 ( .x(n293), .a(dat_o[31]), .b(sel_o[3]) );
    nand2_1 U109 ( .x(n303), .a(dat_o[26]), .b(sel_o[3]) );
    nand2_1 U110 ( .x(n305), .a(dat_o[25]), .b(sel_o[3]) );
    nand2_1 U111 ( .x(n307), .a(dat_o[24]), .b(sel_o[3]) );
    mux2i_1 U113 ( .x(\data[0] ), .d0(n99), .sl(n65), .d1(n222) );
    mux2i_1 U114 ( .x(\data[10] ), .d0(n211), .sl(n214), .d1(n210) );
    mux2i_1 U115 ( .x(\data[11] ), .d0(n209), .sl(n214), .d1(n208) );
    mux2i_1 U116 ( .x(\data[12] ), .d0(n207), .sl(n214), .d1(n206) );
    mux2i_1 U117 ( .x(\data[13] ), .d0(n205), .sl(n214), .d1(n204) );
    mux2i_1 U118 ( .x(\data[14] ), .d0(n63), .sl(n214), .d1(n203) );
    mux2i_1 U119 ( .x(\data[15] ), .d0(n202), .sl(n214), .d1(n201) );
    mux2i_1 U120 ( .x(\data[1] ), .d0(n97), .sl(n65), .d1(n221) );
    mux2i_1 U121 ( .x(\data[2] ), .d0(n95), .sl(n65), .d1(n220) );
    mux2i_1 U122 ( .x(\data[3] ), .d0(n93), .sl(n65), .d1(n219) );
    mux2i_1 U123 ( .x(\data[4] ), .d0(n91), .sl(n65), .d1(n218) );
    mux2i_1 U124 ( .x(\data[5] ), .d0(n89), .sl(n65), .d1(n217) );
    mux2i_1 U125 ( .x(\data[6] ), .d0(n87), .sl(n65), .d1(n216) );
    mux2i_1 U126 ( .x(\data[7] ), .d0(n85), .sl(n65), .d1(n215) );
    mux2i_1 U127 ( .x(\data[8] ), .d0(n200), .sl(n214), .d1(n199) );
    mux2i_1 U128 ( .x(\data[9] ), .d0(n198), .sl(n214), .d1(n197) );
    nor2_1 U129 ( .x(high_ir_rd), .a(n79), .b(n80) );
    mux2i_1 U131 ( .x(\size[0] ), .d0(n212), .sl(n65), .d1(n213) );
    nand2i_1 U132 ( .x(n308), .a(sel_o[1]), .b(n70) );
    inv_1 U133 ( .x(n255), .a(n182) );
    inv_1 U134 ( .x(n256), .a(n179) );
    inv_1 U135 ( .x(n257), .a(n176) );
    inv_1 U136 ( .x(n258), .a(n173) );
    inv_1 U137 ( .x(n260), .a(n194) );
    inv_1 U138 ( .x(n261), .a(n191) );
    inv_1 U139 ( .x(n262), .a(n188) );
    inv_1 U140 ( .x(n263), .a(n185) );
    inv_1 U141 ( .x(n245), .a(n158) );
    inv_1 U142 ( .x(n246), .a(n155) );
    inv_1 U143 ( .x(n247), .a(n152) );
    inv_1 U144 ( .x(n248), .a(n149) );
    inv_1 U145 ( .x(n250), .a(n170) );
    inv_1 U146 ( .x(n251), .a(n167) );
    inv_1 U147 ( .x(n252), .a(n164) );
    inv_1 U148 ( .x(n253), .a(n161) );
    inv_1 U149 ( .x(n235), .a(n134) );
    inv_1 U150 ( .x(n236), .a(n131) );
    inv_1 U151 ( .x(n237), .a(n128) );
    inv_1 U152 ( .x(n238), .a(n125) );
    inv_1 U153 ( .x(n240), .a(n146) );
    inv_1 U154 ( .x(n241), .a(n143) );
    inv_1 U155 ( .x(n242), .a(n140) );
    inv_1 U156 ( .x(n243), .a(n137) );
    inv_1 U157 ( .x(n225), .a(n110) );
    inv_1 U158 ( .x(n226), .a(n107) );
    inv_1 U159 ( .x(n227), .a(n104) );
    inv_1 U160 ( .x(n228), .a(n101) );
    inv_1 U161 ( .x(n230), .a(n122) );
    inv_1 U162 ( .x(n231), .a(n119) );
    inv_1 U163 ( .x(n232), .a(n116) );
    inv_1 U164 ( .x(n233), .a(n113) );
    nor2_1 U165 ( .x(n272), .a(n252), .b(n253) );
    nor2_1 U166 ( .x(n271), .a(n250), .b(n251) );
    nor2_1 U167 ( .x(n275), .a(n247), .b(n248) );
    nor2_1 U168 ( .x(n274), .a(n245), .b(n246) );
    nor2_1 U169 ( .x(n265), .a(n262), .b(n263) );
    nor2_1 U170 ( .x(n264), .a(n260), .b(n261) );
    nor2_1 U171 ( .x(n268), .a(n257), .b(n258) );
    nor2_1 U172 ( .x(n267), .a(n255), .b(n256) );
    nor2_1 U173 ( .x(n286), .a(n232), .b(n233) );
    nor2_1 U174 ( .x(n285), .a(n230), .b(n231) );
    nor2_1 U175 ( .x(n289), .a(n227), .b(n228) );
    nor2_1 U176 ( .x(n288), .a(n225), .b(n226) );
    nor2_1 U177 ( .x(n279), .a(n242), .b(n243) );
    nor2_1 U178 ( .x(n278), .a(n240), .b(n241) );
    nor2_1 U179 ( .x(n282), .a(n237), .b(n238) );
    nor2_1 U180 ( .x(n281), .a(n235), .b(n236) );
    nand2_1 U181 ( .x(n182), .a(n183), .b(n184) );
    nand2_1 U182 ( .x(n179), .a(n180), .b(n181) );
    nand2_1 U183 ( .x(n176), .a(n177), .b(n178) );
    nand2_1 U184 ( .x(n173), .a(n174), .b(n175) );
    nand2_1 U185 ( .x(n194), .a(n195), .b(n196) );
    nand2_1 U186 ( .x(n191), .a(n192), .b(n193) );
    nand2_1 U187 ( .x(n188), .a(n189), .b(n190) );
    nand2_1 U188 ( .x(n185), .a(n186), .b(n187) );
    nand2_1 U189 ( .x(n158), .a(n159), .b(n160) );
    nand2_1 U190 ( .x(n155), .a(n156), .b(n157) );
    nand2_1 U191 ( .x(n152), .a(n153), .b(n154) );
    nand2_1 U192 ( .x(n149), .a(n150), .b(n151) );
    nand2_1 U193 ( .x(n170), .a(n171), .b(n172) );
    nand2_1 U194 ( .x(n167), .a(n168), .b(n169) );
    nand2_1 U195 ( .x(n164), .a(n165), .b(n166) );
    nand2_1 U196 ( .x(n161), .a(n162), .b(n163) );
    nand2_1 U197 ( .x(n134), .a(n135), .b(n136) );
    nand2_1 U198 ( .x(n131), .a(n132), .b(n133) );
    nand2_1 U199 ( .x(n128), .a(n129), .b(n130) );
    nand2_1 U200 ( .x(n125), .a(n126), .b(n127) );
    nand2_1 U201 ( .x(n146), .a(n147), .b(n148) );
    nand2_1 U202 ( .x(n143), .a(n144), .b(n145) );
    nand2_1 U203 ( .x(n140), .a(n141), .b(n142) );
    nand2_1 U204 ( .x(n137), .a(n138), .b(n139) );
    nand2_1 U205 ( .x(n110), .a(n111), .b(n112) );
    nand2_1 U206 ( .x(n107), .a(n108), .b(n109) );
    nand2_1 U207 ( .x(n104), .a(n105), .b(n106) );
    nand2_1 U208 ( .x(n101), .a(n102), .b(n103) );
    nand2_1 U209 ( .x(n122), .a(n123), .b(n124) );
    nand2_1 U210 ( .x(n119), .a(n120), .b(n121) );
    nand2_1 U211 ( .x(n116), .a(n117), .b(n118) );
    nand2_1 U212 ( .x(n113), .a(n114), .b(n115) );
    inv_1 U213 ( .x(n183), .a(ir_rd[60]) );
    inv_1 U214 ( .x(n184), .a(ir_rd[28]) );
    inv_1 U215 ( .x(n180), .a(ir_rd[61]) );
    inv_1 U216 ( .x(n181), .a(ir_rd[29]) );
    inv_1 U217 ( .x(n177), .a(ir_rd[62]) );
    inv_1 U218 ( .x(n178), .a(ir_rd[30]) );
    inv_1 U219 ( .x(n174), .a(ir_rd[63]) );
    inv_1 U220 ( .x(n175), .a(ir_rd[31]) );
    inv_1 U221 ( .x(n195), .a(ir_rd[56]) );
    inv_1 U222 ( .x(n196), .a(ir_rd[24]) );
    inv_1 U223 ( .x(n192), .a(ir_rd[57]) );
    inv_1 U224 ( .x(n193), .a(ir_rd[25]) );
    inv_1 U225 ( .x(n189), .a(ir_rd[58]) );
    inv_1 U226 ( .x(n190), .a(ir_rd[26]) );
    inv_1 U227 ( .x(n186), .a(ir_rd[59]) );
    inv_1 U228 ( .x(n187), .a(ir_rd[27]) );
    inv_1 U229 ( .x(n159), .a(ir_rd[52]) );
    inv_1 U230 ( .x(n160), .a(ir_rd[20]) );
    inv_1 U231 ( .x(n156), .a(ir_rd[53]) );
    inv_1 U232 ( .x(n157), .a(ir_rd[21]) );
    inv_1 U233 ( .x(n153), .a(ir_rd[54]) );
    inv_1 U234 ( .x(n154), .a(ir_rd[22]) );
    inv_1 U235 ( .x(n150), .a(ir_rd[55]) );
    inv_1 U236 ( .x(n151), .a(ir_rd[23]) );
    inv_1 U237 ( .x(n171), .a(ir_rd[48]) );
    inv_1 U238 ( .x(n172), .a(ir_rd[16]) );
    inv_1 U239 ( .x(n168), .a(ir_rd[49]) );
    inv_1 U240 ( .x(n169), .a(ir_rd[17]) );
    inv_1 U241 ( .x(n165), .a(ir_rd[50]) );
    inv_1 U242 ( .x(n166), .a(ir_rd[18]) );
    inv_1 U243 ( .x(n162), .a(ir_rd[51]) );
    inv_1 U244 ( .x(n163), .a(ir_rd[19]) );
    inv_1 U245 ( .x(n135), .a(ir_rd[44]) );
    inv_1 U246 ( .x(n136), .a(ir_rd[12]) );
    inv_1 U247 ( .x(n132), .a(ir_rd[45]) );
    inv_1 U248 ( .x(n133), .a(ir_rd[13]) );
    inv_1 U249 ( .x(n129), .a(ir_rd[46]) );
    inv_1 U250 ( .x(n130), .a(ir_rd[14]) );
    inv_1 U251 ( .x(n126), .a(ir_rd[47]) );
    inv_1 U252 ( .x(n127), .a(ir_rd[15]) );
    inv_1 U253 ( .x(n147), .a(ir_rd[40]) );
    inv_1 U254 ( .x(n148), .a(ir_rd[8]) );
    inv_1 U255 ( .x(n144), .a(ir_rd[41]) );
    inv_1 U256 ( .x(n145), .a(ir_rd[9]) );
    inv_1 U257 ( .x(n141), .a(ir_rd[42]) );
    inv_1 U258 ( .x(n142), .a(ir_rd[10]) );
    inv_1 U259 ( .x(n138), .a(ir_rd[43]) );
    inv_1 U260 ( .x(n139), .a(ir_rd[11]) );
    inv_1 U261 ( .x(n111), .a(ir_rd[36]) );
    inv_1 U262 ( .x(n108), .a(ir_rd[37]) );
    inv_1 U263 ( .x(n109), .a(ir_rd[5]) );
    inv_1 U264 ( .x(n105), .a(ir_rd[38]) );
    inv_1 U265 ( .x(n106), .a(ir_rd[6]) );
    inv_1 U266 ( .x(n102), .a(ir_rd[39]) );
    inv_1 U267 ( .x(n103), .a(ir_rd[7]) );
    inv_1 U268 ( .x(n123), .a(ir_rd[32]) );
    inv_1 U269 ( .x(n120), .a(ir_rd[33]) );
    inv_1 U270 ( .x(n121), .a(ir_rd[1]) );
    inv_1 U271 ( .x(n117), .a(ir_rd[34]) );
    inv_1 U272 ( .x(n114), .a(ir_rd[35]) );
    inv_1 U273 ( .x(n115), .a(ir_rd[3]) );
    latn_1 \dat_i_reg[30]  ( .q(dat_i[30]), .d(ir_rd[62]), .g(n7) );
    latn_1 \dat_i_reg[28]  ( .q(dat_i[28]), .d(ir_rd[60]), .g(n7) );
    latn_1 \dat_i_reg[27]  ( .q(dat_i[27]), .d(ir_rd[59]), .g(n7) );
    latn_1 \dat_i_reg[26]  ( .q(dat_i[26]), .d(ir_rd[58]), .g(n7) );
    latn_1 \dat_i_reg[25]  ( .q(dat_i[25]), .d(ir_rd[57]), .g(n7) );
    latn_1 \dat_i_reg[24]  ( .q(dat_i[24]), .d(ir_rd[56]), .g(n7) );
    latn_1 \dat_i_reg[22]  ( .q(dat_i[22]), .d(ir_rd[54]), .g(n7) );
    latn_1 \dat_i_reg[20]  ( .q(dat_i[20]), .d(ir_rd[52]), .g(n7) );
    latn_1 \dat_i_reg[19]  ( .q(dat_i[19]), .d(ir_rd[51]), .g(n7) );
    latn_1 \dat_i_reg[18]  ( .q(dat_i[18]), .d(ir_rd[50]), .g(n7) );
    latn_1 \dat_i_reg[17]  ( .q(dat_i[17]), .d(ir_rd[49]), .g(n7) );
    latn_1 \dat_i_reg[16]  ( .q(dat_i[16]), .d(ir_rd[48]), .g(n6) );
    latn_1 \dat_i_reg[14]  ( .q(dat_i[14]), .d(ir_rd[46]), .g(n6) );
    latn_1 \dat_i_reg[12]  ( .q(dat_i[12]), .d(ir_rd[44]), .g(n6) );
    latn_1 \dat_i_reg[10]  ( .q(dat_i[10]), .d(ir_rd[42]), .g(n6) );
    latn_1 \dat_i_reg[8]  ( .q(dat_i[8]), .d(ir_rd[40]), .g(n6) );
    latn_1 \dat_i_reg[6]  ( .q(dat_i[6]), .d(ir_rd[38]), .g(n6) );
    latn_1 \dat_i_reg[4]  ( .q(dat_i[4]), .d(ir_rd[36]), .g(n6) );
    latn_1 \dat_i_reg[3]  ( .q(dat_i[3]), .d(ir_rd[35]), .g(n1) );
    latn_1 \dat_i_reg[2]  ( .q(dat_i[2]), .d(ir_rd[34]), .g(n1) );
    latn_1 \dat_i_reg[1]  ( .q(dat_i[1]), .d(ir_rd[33]), .g(n1) );
    latn_1 \dat_i_reg[0]  ( .q(dat_i[0]), .d(ir_rd[32]), .g(n1) );
    latn_1 we_i_reg ( .q(we_i), .d(ir_rnw[0]), .g(n1) );
    latn_1 err_i_reg ( .q(err_i), .d(ir_err[1]), .g(n1) );
    latn_1 \dat_i_reg[13]  ( .q(dat_i[13]), .d(ir_rd[45]), .g(n6) );
    latn_1 \dat_i_reg[5]  ( .q(dat_i[5]), .d(ir_rd[37]), .g(n1) );
    latn_1 \dat_i_reg[15]  ( .q(dat_i[15]), .d(ir_rd[47]), .g(n6) );
    latn_1 \dat_i_reg[7]  ( .q(dat_i[7]), .d(ir_rd[39]), .g(n1) );
    latn_1 \dat_i_reg[29]  ( .q(dat_i[29]), .d(ir_rd[61]), .g(n6) );
    latn_1 \dat_i_reg[21]  ( .q(dat_i[21]), .d(ir_rd[53]), .g(n1) );
    latn_1 \dat_i_reg[31]  ( .q(dat_i[31]), .d(ir_rd[63]), .g(n6) );
    latn_1 \dat_i_reg[23]  ( .q(dat_i[23]), .d(ir_rd[55]), .g(n1) );
    latn_1 \dat_i_reg[9]  ( .q(dat_i[9]), .d(ir_rd[41]), .g(n6) );
    latn_1 \dat_i_reg[11]  ( .q(dat_i[11]), .d(ir_rd[43]), .g(n1) );
    oa21_1 \all_write/__tmp99/U1  ( .x(all_w), .a(_28_net_), .b(all_w), .c(
        comp_basic) );
    ao31_1 \all_read/__tmp99/aoi  ( .x(\all_read/__tmp99/loop ), .a(comp_basic
        ), .b(comp_rd), .c(_27_net_), .d(all_r) );
    oa21_1 \all_read/__tmp99/outGate  ( .x(all_r), .a(comp_basic), .b(comp_rd), 
        .c(\all_read/__tmp99/loop ) );
    ao222_1 \rd/__tmp99/U1  ( .x(comp_rd), .a(high_ir_rd), .b(low_ir_rd), .c(
        high_ir_rd), .d(comp_rd), .e(low_ir_rd), .f(comp_rd) );
    ao222_1 \basic/__tmp99/U1  ( .x(comp_basic), .a(_25_net_), .b(_26_net_), 
        .c(_25_net_), .d(comp_basic), .e(_26_net_), .f(comp_basic) );
    inv_1 \Ucol2/Uii  ( .x(\Ucol2/ni ), .a(ts_o[2]) );
    inv_1 \Ucol2/Uih  ( .x(\Ucol2/nh ), .a(ic_col[5]) );
    inv_1 \Ucol2/Uil  ( .x(\Ucol2/nl ), .a(ic_col[2]) );
    ao23_1 \Ucol2/Ucl/U1/U1  ( .x(ic_col[2]), .a(n11), .b(ic_col[2]), .c(n8), 
        .d(\Ucol2/ni ), .e(\Ucol2/nh ) );
    ao23_1 \Ucol2/Uch/U1/U1  ( .x(ic_col[5]), .a(n11), .b(ic_col[5]), .c(n8), 
        .d(ts_o[2]), .e(\Ucol2/nl ) );
    inv_1 \Ucol1/Uii  ( .x(\Ucol1/ni ), .a(ts_o[1]) );
    inv_1 \Ucol1/Uih  ( .x(\Ucol1/nh ), .a(ic_col[4]) );
    inv_1 \Ucol1/Uil  ( .x(\Ucol1/nl ), .a(ic_col[1]) );
    ao23_1 \Ucol1/Ucl/U1/U1  ( .x(ic_col[1]), .a(n11), .b(ic_col[1]), .c(n8), 
        .d(\Ucol1/ni ), .e(\Ucol1/nh ) );
    ao23_1 \Ucol1/Uch/U1/U1  ( .x(ic_col[4]), .a(n11), .b(ic_col[4]), .c(n9), 
        .d(ts_o[1]), .e(\Ucol1/nl ) );
    inv_1 \Ucol0/Uii  ( .x(\Ucol0/ni ), .a(ts_o[0]) );
    inv_1 \Ucol0/Uih  ( .x(\Ucol0/nh ), .a(ic_col[3]) );
    inv_1 \Ucol0/Uil  ( .x(\Ucol0/nl ), .a(ic_col[0]) );
    ao23_1 \Ucol0/Ucl/U1/U1  ( .x(ic_col[0]), .a(n11), .b(ic_col[0]), .c(n10), 
        .d(\Ucol0/ni ), .e(\Ucol0/nh ) );
    ao23_1 \Ucol0/Uch/U1/U1  ( .x(ic_col[3]), .a(n11), .b(ic_col[3]), .c(n9), 
        .d(ts_o[0]), .e(\Ucol0/nl ) );
    inv_1 \Utag4/Uii  ( .x(\Utag4/ni ), .a(tag_id[4]) );
    inv_1 \Utag4/Uih  ( .x(\Utag4/nh ), .a(ic_itag[9]) );
    inv_1 \Utag4/Uil  ( .x(\Utag4/nl ), .a(ic_itag[4]) );
    ao23_1 \Utag4/Ucl/U1/U1  ( .x(ic_itag[4]), .a(n11), .b(ic_itag[4]), .c(n9), 
        .d(\Utag4/ni ), .e(\Utag4/nh ) );
    ao23_1 \Utag4/Uch/U1/U1  ( .x(ic_itag[9]), .a(n10), .b(ic_itag[9]), .c(n9), 
        .d(tag_id[4]), .e(\Utag4/nl ) );
    inv_1 \Utag3/Uii  ( .x(\Utag3/ni ), .a(tag_id[3]) );
    inv_1 \Utag3/Uih  ( .x(\Utag3/nh ), .a(ic_itag[8]) );
    inv_1 \Utag3/Uil  ( .x(\Utag3/nl ), .a(ic_itag[3]) );
    ao23_1 \Utag3/Ucl/U1/U1  ( .x(ic_itag[3]), .a(n10), .b(ic_itag[3]), .c(n9), 
        .d(\Utag3/ni ), .e(\Utag3/nh ) );
    ao23_1 \Utag3/Uch/U1/U1  ( .x(ic_itag[8]), .a(n10), .b(ic_itag[8]), .c(n9), 
        .d(tag_id[3]), .e(\Utag3/nl ) );
    inv_1 \Utag2/Uii  ( .x(\Utag2/ni ), .a(tag_id[2]) );
    inv_1 \Utag2/Uih  ( .x(\Utag2/nh ), .a(ic_itag[7]) );
    inv_1 \Utag2/Uil  ( .x(\Utag2/nl ), .a(ic_itag[2]) );
    ao23_1 \Utag2/Ucl/U1/U1  ( .x(ic_itag[2]), .a(n10), .b(ic_itag[2]), .c(n9), 
        .d(\Utag2/ni ), .e(\Utag2/nh ) );
    ao23_1 \Utag2/Uch/U1/U1  ( .x(ic_itag[7]), .a(n10), .b(ic_itag[7]), .c(n10
        ), .d(tag_id[2]), .e(\Utag2/nl ) );
    inv_1 \Utag1/Uii  ( .x(\Utag1/ni ), .a(tag_id[1]) );
    inv_1 \Utag1/Uih  ( .x(\Utag1/nh ), .a(ic_itag[6]) );
    inv_1 \Utag1/Uil  ( .x(\Utag1/nl ), .a(ic_itag[1]) );
    ao23_1 \Utag1/Ucl/U1/U1  ( .x(ic_itag[1]), .a(n11), .b(ic_itag[1]), .c(n9), 
        .d(\Utag1/ni ), .e(\Utag1/nh ) );
    ao23_1 \Utag1/Uch/U1/U1  ( .x(ic_itag[6]), .a(n11), .b(ic_itag[6]), .c(n9), 
        .d(tag_id[1]), .e(\Utag1/nl ) );
    inv_1 \Utag0/Uii  ( .x(\Utag0/ni ), .a(tag_id[0]) );
    inv_1 \Utag0/Uih  ( .x(\Utag0/nh ), .a(ic_itag[5]) );
    inv_1 \Utag0/Uil  ( .x(\Utag0/nl ), .a(ic_itag[0]) );
    ao23_1 \Utag0/Ucl/U1/U1  ( .x(ic_itag[0]), .a(n11), .b(ic_itag[0]), .c(n8), 
        .d(\Utag0/ni ), .e(\Utag0/nh ) );
    ao23_1 \Utag0/Uch/U1/U1  ( .x(ic_itag[5]), .a(n10), .b(ic_itag[5]), .c(n8), 
        .d(tag_id[0]), .e(\Utag0/nl ) );
    inv_1 \Usze1/Uii  ( .x(\Usze1/ni ), .a(\size[1] ) );
    inv_1 \Usze1/Uih  ( .x(\Usze1/nh ), .a(ic_size[3]) );
    inv_1 \Usze1/Uil  ( .x(\Usze1/nl ), .a(ic_size[1]) );
    ao23_1 \Usze1/Ucl/U1/U1  ( .x(ic_size[1]), .a(n10), .b(ic_size[1]), .c(n9), 
        .d(\Usze1/ni ), .e(\Usze1/nh ) );
    ao23_1 \Usze1/Uch/U1/U1  ( .x(ic_size[3]), .a(n10), .b(ic_size[3]), .c(n9), 
        .d(\size[1] ), .e(\Usze1/nl ) );
    inv_1 \Usze0/Uii  ( .x(\Usze0/ni ), .a(\size[0] ) );
    inv_1 \Usze0/Uih  ( .x(\Usze0/nh ), .a(ic_size[2]) );
    inv_1 \Usze0/Uil  ( .x(\Usze0/nl ), .a(ic_size[0]) );
    ao23_1 \Usze0/Ucl/U1/U1  ( .x(ic_size[0]), .a(n10), .b(ic_size[0]), .c(n9), 
        .d(\Usze0/ni ), .e(\Usze0/nh ) );
    ao23_1 \Usze0/Uch/U1/U1  ( .x(ic_size[2]), .a(n10), .b(ic_size[2]), .c(n9), 
        .d(\size[0] ), .e(\Usze0/nl ) );
    inv_1 \Urnw/Uii  ( .x(\Urnw/ni ), .a(_24_net_) );
    inv_1 \Urnw/Uih  ( .x(\Urnw/nh ), .a(ic_rnw[1]) );
    inv_1 \Urnw/Uil  ( .x(\Urnw/nl ), .a(ic_rnw[0]) );
    ao23_1 \Urnw/Ucl/U1/U1  ( .x(ic_rnw[0]), .a(n10), .b(ic_rnw[0]), .c(n9), 
        .d(\Urnw/ni ), .e(\Urnw/nh ) );
    ao23_1 \Urnw/Uch/U1/U1  ( .x(ic_rnw[1]), .a(n10), .b(ic_rnw[1]), .c(n9), 
        .d(_24_net_), .e(\Urnw/nl ) );
    inv_1 \Ulock/Uii  ( .x(\Ulock/ni ), .a(mult_o) );
    inv_1 \Ulock/Uih  ( .x(\Ulock/nh ), .a(ic_lock[1]) );
    inv_1 \Ulock/Uil  ( .x(\Ulock/nl ), .a(ic_lock[0]) );
    ao23_1 \Ulock/Ucl/U1/U1  ( .x(ic_lock[0]), .a(n11), .b(ic_lock[0]), .c(n9), 
        .d(\Ulock/ni ), .e(\Ulock/nh ) );
    ao23_1 \Ulock/Uch/U1/U1  ( .x(ic_lock[1]), .a(n11), .b(ic_lock[1]), .c(n8), 
        .d(mult_o), .e(\Ulock/nl ) );
    inv_1 \Upred/Uii  ( .x(\Upred/ni ), .a(prd_o) );
    inv_1 \Upred/Uih  ( .x(\Upred/nh ), .a(ic_pred[1]) );
    inv_1 \Upred/Uil  ( .x(\Upred/nl ), .a(ic_pred[0]) );
    ao23_1 \Upred/Ucl/U1/U1  ( .x(ic_pred[0]), .a(n11), .b(ic_pred[0]), .c(n8), 
        .d(\Upred/ni ), .e(\Upred/nh ) );
    ao23_1 \Upred/Uch/U1/U1  ( .x(ic_pred[1]), .a(n10), .b(ic_pred[1]), .c(n8), 
        .d(prd_o), .e(\Upred/nl ) );
    inv_1 \Useq/Uii  ( .x(\Useq/ni ), .a(seq_o) );
    inv_1 \Useq/Uih  ( .x(\Useq/nh ), .a(ic_seq[1]) );
    inv_1 \Useq/Uil  ( .x(\Useq/nl ), .a(ic_seq[0]) );
    ao23_1 \Useq/Ucl/U1/U1  ( .x(ic_seq[0]), .a(n10), .b(ic_seq[0]), .c(n8), 
        .d(\Useq/ni ), .e(\Useq/nh ) );
    ao23_1 \Useq/Uch/U1/U1  ( .x(ic_seq[1]), .a(n11), .b(ic_seq[1]), .c(n8), 
        .d(seq_o), .e(\Useq/nl ) );
    buf_3 U1 ( .x(n1), .a(en) );
    buf_3 U41 ( .x(n7), .a(en) );
    buf_3 U43 ( .x(n6), .a(en) );
    inv_2 U44 ( .x(n214), .a(n308) );
    buf_3 U47 ( .x(n65), .a(sel_o[0]) );
    nand3i_0 U49 ( .x(n212), .a(sel_o[1]), .b(sel_o[3]), .c(n70) );
    nor2_0 U50 ( .x(n223), .a(n70), .b(sel_o[3]) );
    nand2_0 U58 ( .x(n297), .a(dat_o[29]), .b(sel_o[3]) );
    nand2_0 U102 ( .x(n301), .a(dat_o[27]), .b(sel_o[3]) );
    nand2_0 U105 ( .x(n299), .a(dat_o[28]), .b(sel_o[3]) );
    nand2_0 U106 ( .x(n295), .a(dat_o[30]), .b(sel_o[3]) );
    inv_0 U107 ( .x(n78), .a(ir_err[0]) );
    buf_16 U108 ( .x(n8), .a(req_in_delayed) );
    buf_16 U279 ( .x(n9), .a(req_in_delayed) );
    buf_16 U280 ( .x(n10), .a(req_in_delayed) );
    buf_16 U281 ( .x(n11), .a(req_in_delayed) );
endmodule


module master_if_dport ( nReset, mc_req, mc_we, mc_mult, mc_prd, mc_seq, mc_ts, 
    mc_sel, mc_adr, mc_dat, mc_ack, mr_req, mr_we, mr_err, mr_rty, mr_acc, 
    mr_ts, mr_sel, mr_dat, mr_ack, chaincommand, nchaincommandack, 
    chainresponse, nchainresponseack, e_bare, e_dm, e_im, e_wish, r_bare, r_dm, 
    r_im, r_wish, tag_id, force_bare );
input  [2:0] mc_ts;
input  [3:0] mc_sel;
input  [31:0] mc_adr;
input  [31:0] mc_dat;
output [2:0] mr_ts;
output [3:0] mr_sel;
output [31:0] mr_dat;
output [4:0] chaincommand;
input  [4:0] chainresponse;
input  [3:0] e_bare;
input  [3:0] e_dm;
input  [3:0] e_im;
input  [3:0] e_wish;
input  [3:0] r_bare;
input  [3:0] r_dm;
input  [3:0] r_im;
input  [3:0] r_wish;
input  [4:0] tag_id;
input  nReset, mc_req, mc_we, mc_mult, mc_prd, mc_seq, mr_ack, 
    nchaincommandack, force_bare;
output mc_ack, mr_req, mr_we, mr_err, mr_rty, mr_acc, nchainresponseack;
    wire \ci_seq[1] , \ci_seq[0] , \ci_lock[1] , \ci_lock[0] , \ci_rnw[1] , 
        \ci_rnw[0] , \ci_size[3] , \ci_size[2] , \ci_size[1] , \ci_size[0] , 
        \ci_itag[9] , \ci_itag[8] , \ci_itag[7] , \ci_itag[6] , \ci_itag[5] , 
        \ci_itag[4] , \ci_itag[3] , \ci_itag[2] , \ci_itag[1] , \ci_itag[0] , 
        \ci_a[63] , \ci_a[62] , \ci_a[61] , \ci_a[60] , \ci_a[59] , \ci_a[58] , 
        \ci_a[57] , \ci_a[56] , \ci_a[55] , \ci_a[54] , \ci_a[53] , \ci_a[52] , 
        \ci_a[51] , \ci_a[50] , \ci_a[49] , \ci_a[48] , \ci_a[47] , \ci_a[46] , 
        \ci_a[45] , \ci_a[44] , \ci_a[43] , \ci_a[42] , \ci_a[41] , \ci_a[40] , 
        \ci_a[39] , \ci_a[38] , \ci_a[37] , \ci_a[36] , \ci_a[35] , \ci_a[34] , 
        \ci_a[33] , \ci_a[32] , \ci_a[31] , \ci_a[30] , \ci_a[29] , \ci_a[28] , 
        \ci_a[27] , \ci_a[26] , \ci_a[25] , \ci_a[24] , \ci_a[23] , \ci_a[22] , 
        \ci_a[21] , \ci_a[20] , \ci_a[19] , \ci_a[18] , \ci_a[17] , \ci_a[16] , 
        \ci_a[15] , \ci_a[14] , \ci_a[13] , \ci_a[12] , \ci_a[11] , \ci_a[10] , 
        \ci_a[9] , \ci_a[8] , \ci_a[7] , \ci_a[6] , \ci_a[5] , \ci_a[4] , 
        \ci_a[3] , \ci_a[2] , \ci_a[1] , \ci_a[0] , \ci_wd[63] , \ci_wd[62] , 
        \ci_wd[61] , \ci_wd[60] , \ci_wd[59] , \ci_wd[58] , \ci_wd[57] , 
        \ci_wd[56] , \ci_wd[55] , \ci_wd[54] , \ci_wd[53] , \ci_wd[52] , 
        \ci_wd[51] , \ci_wd[50] , \ci_wd[49] , \ci_wd[48] , \ci_wd[47] , 
        \ci_wd[46] , \ci_wd[45] , \ci_wd[44] , \ci_wd[43] , \ci_wd[42] , 
        \ci_wd[41] , \ci_wd[40] , \ci_wd[39] , \ci_wd[38] , \ci_wd[37] , 
        \ci_wd[36] , \ci_wd[35] , \ci_wd[34] , \ci_wd[33] , \ci_wd[32] , 
        \ci_wd[31] , \ci_wd[30] , \ci_wd[29] , \ci_wd[28] , \ci_wd[27] , 
        \ci_wd[26] , \ci_wd[25] , \ci_wd[24] , \ci_wd[23] , \ci_wd[22] , 
        \ci_wd[21] , \ci_wd[20] , \ci_wd[19] , \ci_wd[18] , \ci_wd[17] , 
        \ci_wd[16] , \ci_wd[15] , \ci_wd[14] , \ci_wd[13] , \ci_wd[12] , 
        \ci_wd[11] , \ci_wd[10] , \ci_wd[9] , \ci_wd[8] , \ci_wd[7] , 
        \ci_wd[6] , \ci_wd[5] , \ci_wd[4] , \ci_wd[3] , \ci_wd[2] , \ci_wd[1] , 
        \ci_wd[0] , \ci_pred[1] , \ci_pred[0] , \ci_col[5] , \ci_col[4] , 
        \ci_col[3] , \ci_col[2] , \ci_col[1] , \ci_col[0] , ci_ack, 
        \ri_err[1] , \ri_err[0] , \ri_rnw[1] , \ri_rnw[0] , \ri_rd[63] , 
        \ri_rd[62] , \ri_rd[61] , \ri_rd[60] , \ri_rd[59] , \ri_rd[58] , 
        \ri_rd[57] , \ri_rd[56] , \ri_rd[55] , \ri_rd[54] , \ri_rd[53] , 
        \ri_rd[52] , \ri_rd[51] , \ri_rd[50] , \ri_rd[49] , \ri_rd[48] , 
        \ri_rd[47] , \ri_rd[46] , \ri_rd[45] , \ri_rd[44] , \ri_rd[43] , 
        \ri_rd[42] , \ri_rd[41] , \ri_rd[40] , \ri_rd[39] , \ri_rd[38] , 
        \ri_rd[37] , \ri_rd[36] , \ri_rd[35] , \ri_rd[34] , \ri_rd[33] , 
        \ri_rd[32] , \ri_rd[31] , \ri_rd[30] , \ri_rd[29] , \ri_rd[28] , 
        \ri_rd[27] , \ri_rd[26] , \ri_rd[25] , \ri_rd[24] , \ri_rd[23] , 
        \ri_rd[22] , \ri_rd[21] , \ri_rd[20] , \ri_rd[19] , \ri_rd[18] , 
        \ri_rd[17] , \ri_rd[16] , \ri_rd[15] , \ri_rd[14] , \ri_rd[13] , 
        \ri_rd[12] , \ri_rd[11] , \ri_rd[10] , \ri_rd[9] , \ri_rd[8] , 
        \ri_rd[7] , \ri_rd[6] , \ri_rd[5] , \ri_rd[4] , \ri_rd[3] , \ri_rd[2] , 
        \ri_rd[1] , \ri_rd[0] , ri_ack, reset, nroute_ack, routetx_req, 
        routetx_ack, \route[4] , \route[1] , \route[0] , \i_eh[2] , \i_eh[1] , 
        \i_eh[0] , \i_el[3] , \i_el[2] , \i_el[1] , \i_el[0] , \i_rh[3] , 
        \i_rh[2] , \i_rh[1] , \i_rl[3] , \i_rl[2] , \i_rl[1] , \i_rl[0] ;
    wire SYNOPSYS_UNCONNECTED_1 , SYNOPSYS_UNCONNECTED_2 , 
	SYNOPSYS_UNCONNECTED_3 , SYNOPSYS_UNCONNECTED_4 ;
    assign mr_rty = 1'b0;
    assign mr_acc = 1'b0;
    assign mr_ts[2] = 1'b0;
    assign mr_ts[1] = 1'b0;
    assign mr_ts[0] = 1'b0;
    assign mr_sel[3] = 1'b0;
    assign mr_sel[2] = 1'b0;
    assign mr_sel[1] = 1'b0;
    assign mr_sel[0] = 1'b0;
    inv_2 U1 ( .x(reset), .a(nReset) );
    m2cp_dport master2chainif ( .req_in(mc_req), .ts_o(mc_ts), .sel_o(mc_sel), 
        .mult_o(mc_mult), .we_o(mc_we), .prd_o(mc_prd), .seq_o(mc_seq), 
        .adr_o(mc_adr), .dat_o(mc_dat), .ain(mc_ack), .ic_seq({\ci_seq[1] , 
        \ci_seq[0] }), .ic_pred({\ci_pred[1] , \ci_pred[0] }), .ic_size({
        \ci_size[3] , \ci_size[2] , \ci_size[1] , \ci_size[0] }), .ic_itag({
        \ci_itag[9] , \ci_itag[8] , \ci_itag[7] , \ci_itag[6] , \ci_itag[5] , 
        \ci_itag[4] , \ci_itag[3] , \ci_itag[2] , \ci_itag[1] , \ci_itag[0] }), 
        .ic_wd({\ci_wd[63] , \ci_wd[62] , \ci_wd[61] , \ci_wd[60] , 
        \ci_wd[59] , \ci_wd[58] , \ci_wd[57] , \ci_wd[56] , \ci_wd[55] , 
        \ci_wd[54] , \ci_wd[53] , \ci_wd[52] , \ci_wd[51] , \ci_wd[50] , 
        \ci_wd[49] , \ci_wd[48] , \ci_wd[47] , \ci_wd[46] , \ci_wd[45] , 
        \ci_wd[44] , \ci_wd[43] , \ci_wd[42] , \ci_wd[41] , \ci_wd[40] , 
        \ci_wd[39] , \ci_wd[38] , \ci_wd[37] , \ci_wd[36] , \ci_wd[35] , 
        \ci_wd[34] , \ci_wd[33] , \ci_wd[32] , \ci_wd[31] , \ci_wd[30] , 
        \ci_wd[29] , \ci_wd[28] , \ci_wd[27] , \ci_wd[26] , \ci_wd[25] , 
        \ci_wd[24] , \ci_wd[23] , \ci_wd[22] , \ci_wd[21] , \ci_wd[20] , 
        \ci_wd[19] , \ci_wd[18] , \ci_wd[17] , \ci_wd[16] , \ci_wd[15] , 
        \ci_wd[14] , \ci_wd[13] , \ci_wd[12] , \ci_wd[11] , \ci_wd[10] , 
        \ci_wd[9] , \ci_wd[8] , \ci_wd[7] , \ci_wd[6] , \ci_wd[5] , \ci_wd[4] , 
        \ci_wd[3] , \ci_wd[2] , \ci_wd[1] , \ci_wd[0] }), .ic_lock({
        \ci_lock[1] , \ci_lock[0] }), .ic_a({\ci_a[63] , \ci_a[62] , 
        \ci_a[61] , \ci_a[60] , \ci_a[59] , \ci_a[58] , \ci_a[57] , \ci_a[56] , 
        \ci_a[55] , \ci_a[54] , \ci_a[53] , \ci_a[52] , \ci_a[51] , \ci_a[50] , 
        \ci_a[49] , \ci_a[48] , \ci_a[47] , \ci_a[46] , \ci_a[45] , \ci_a[44] , 
        \ci_a[43] , \ci_a[42] , \ci_a[41] , \ci_a[40] , \ci_a[39] , \ci_a[38] , 
        \ci_a[37] , \ci_a[36] , \ci_a[35] , \ci_a[34] , \ci_a[33] , \ci_a[32] , 
        \ci_a[31] , \ci_a[30] , \ci_a[29] , \ci_a[28] , \ci_a[27] , \ci_a[26] , 
        \ci_a[25] , \ci_a[24] , \ci_a[23] , \ci_a[22] , \ci_a[21] , \ci_a[20] , 
        \ci_a[19] , \ci_a[18] , \ci_a[17] , \ci_a[16] , \ci_a[15] , \ci_a[14] , 
        \ci_a[13] , \ci_a[12] , \ci_a[11] , \ci_a[10] , \ci_a[9] , \ci_a[8] , 
        \ci_a[7] , \ci_a[6] , \ci_a[5] , \ci_a[4] , \ci_a[3] , \ci_a[2] , 
        \ci_a[1] , \ci_a[0] }), .ic_rnw({\ci_rnw[1] , \ci_rnw[0] }), .ic_col({
        \ci_col[5] , \ci_col[4] , \ci_col[3] , \ci_col[2] , \ci_col[1] , 
        \ci_col[0] }), .ic_ack(ci_ack), .req_out(mr_req), .we_i(mr_we), 
        .err_i(mr_err), .dat_i(mr_dat), .aout(mr_ack), .ir_rd({\ri_rd[63] , 
        \ri_rd[62] , \ri_rd[61] , \ri_rd[60] , \ri_rd[59] , \ri_rd[58] , 
        \ri_rd[57] , \ri_rd[56] , \ri_rd[55] , \ri_rd[54] , \ri_rd[53] , 
        \ri_rd[52] , \ri_rd[51] , \ri_rd[50] , \ri_rd[49] , \ri_rd[48] , 
        \ri_rd[47] , \ri_rd[46] , \ri_rd[45] , \ri_rd[44] , \ri_rd[43] , 
        \ri_rd[42] , \ri_rd[41] , \ri_rd[40] , \ri_rd[39] , \ri_rd[38] , 
        \ri_rd[37] , \ri_rd[36] , \ri_rd[35] , \ri_rd[34] , \ri_rd[33] , 
        \ri_rd[32] , \ri_rd[31] , \ri_rd[30] , \ri_rd[29] , \ri_rd[28] , 
        \ri_rd[27] , \ri_rd[26] , \ri_rd[25] , \ri_rd[24] , \ri_rd[23] , 
        \ri_rd[22] , \ri_rd[21] , \ri_rd[20] , \ri_rd[19] , \ri_rd[18] , 
        \ri_rd[17] , \ri_rd[16] , \ri_rd[15] , \ri_rd[14] , \ri_rd[13] , 
        \ri_rd[12] , \ri_rd[11] , \ri_rd[10] , \ri_rd[9] , \ri_rd[8] , 
        \ri_rd[7] , \ri_rd[6] , \ri_rd[5] , \ri_rd[4] , \ri_rd[3] , \ri_rd[2] , 
        \ri_rd[1] , \ri_rd[0] }), .ir_err({\ri_err[1] , \ri_err[0] }), 
        .ir_rnw({\ri_rnw[1] , \ri_rnw[0] }), .ir_ack(ri_ack), .tag_id(tag_id), 
        .reset(reset) );
    i_adec_dport dec ( .e_h({SYNOPSYS_UNCONNECTED_1, \i_eh[2] , \i_eh[1] , 
        \i_eh[0] }), .e_l({\i_el[3] , \i_el[2] , \i_el[1] , \i_el[0] }), .r_h(
        {\i_rh[3] , \i_rh[2] , \i_rh[1] , SYNOPSYS_UNCONNECTED_2}), .r_l({
        \i_rl[3] , \i_rl[2] , \i_rl[1] , \i_rl[0] }), .ah({\ci_a[63] , 
        \ci_a[62] , \ci_a[61] , \ci_a[60] , \ci_a[59] , \ci_a[58] , \ci_a[57] , 
        \ci_a[56] , \ci_a[55] , \ci_a[54] , \ci_a[53] , \ci_a[52] , \ci_a[51] , 
        \ci_a[50] , \ci_a[49] , \ci_a[48] , \ci_a[47] , \ci_a[46] , \ci_a[45] , 
        \ci_a[44] , \ci_a[43] , \ci_a[42] , \ci_a[41] , \ci_a[40] , \ci_a[39] , 
        \ci_a[38] , \ci_a[37] , \ci_a[36] , \ci_a[35] , \ci_a[34] , \ci_a[33] , 
        \ci_a[32] }), .al({\ci_a[31] , \ci_a[30] , \ci_a[29] , \ci_a[28] , 
        \ci_a[27] , \ci_a[26] , \ci_a[25] , \ci_a[24] , \ci_a[23] , \ci_a[22] , 
        \ci_a[21] , \ci_a[20] , \ci_a[19] , \ci_a[18] , \ci_a[17] , \ci_a[16] , 
        \ci_a[15] , \ci_a[14] , \ci_a[13] , \ci_a[12] , \ci_a[11] , \ci_a[10] , 
        \ci_a[9] , \ci_a[8] , \ci_a[7] , \ci_a[6] , \ci_a[5] , \ci_a[4] , 
        \ci_a[3] , \ci_a[2] , \ci_a[1] , \ci_a[0] }), .e_bare(e_bare), .e_dm(
        e_dm), .e_im(e_im), .e_wish(e_wish), .r_bare(r_bare), .r_dm(r_dm), 
        .r_im(r_im), .r_wish(r_wish), .force_bare(force_bare) );
    route_tx_dport rt ( .o({\route[4] , SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, \route[1] , \route[0] }), .rtxack(routetx_ack), 
        .e_h({1'b0, \i_eh[2] , \i_eh[1] , \i_eh[0] }), .e_l({\i_el[3] , 
        \i_el[2] , \i_el[1] , \i_el[0] }), .noa(nroute_ack), .r_h({\i_rh[3] , 
        \i_rh[2] , \i_rh[1] , 1'b0}), .r_l({\i_rl[3] , \i_rl[2] , \i_rl[1] , 
        \i_rl[0] }), .rtxreq(routetx_req) );
    initiator_dport it ( .cack(ci_ack), .chaincommand(chaincommand), .err({
        \ri_err[1] , \ri_err[0] }), .nchainresponseack(nchainresponseack), 
        .nrouteack(nroute_ack), .rd({\ri_rd[63] , \ri_rd[62] , \ri_rd[61] , 
        \ri_rd[60] , \ri_rd[59] , \ri_rd[58] , \ri_rd[57] , \ri_rd[56] , 
        \ri_rd[55] , \ri_rd[54] , \ri_rd[53] , \ri_rd[52] , \ri_rd[51] , 
        \ri_rd[50] , \ri_rd[49] , \ri_rd[48] , \ri_rd[47] , \ri_rd[46] , 
        \ri_rd[45] , \ri_rd[44] , \ri_rd[43] , \ri_rd[42] , \ri_rd[41] , 
        \ri_rd[40] , \ri_rd[39] , \ri_rd[38] , \ri_rd[37] , \ri_rd[36] , 
        \ri_rd[35] , \ri_rd[34] , \ri_rd[33] , \ri_rd[32] , \ri_rd[31] , 
        \ri_rd[30] , \ri_rd[29] , \ri_rd[28] , \ri_rd[27] , \ri_rd[26] , 
        \ri_rd[25] , \ri_rd[24] , \ri_rd[23] , \ri_rd[22] , \ri_rd[21] , 
        \ri_rd[20] , \ri_rd[19] , \ri_rd[18] , \ri_rd[17] , \ri_rd[16] , 
        \ri_rd[15] , \ri_rd[14] , \ri_rd[13] , \ri_rd[12] , \ri_rd[11] , 
        \ri_rd[10] , \ri_rd[9] , \ri_rd[8] , \ri_rd[7] , \ri_rd[6] , 
        \ri_rd[5] , \ri_rd[4] , \ri_rd[3] , \ri_rd[2] , \ri_rd[1] , \ri_rd[0] 
        }), .routetxreq(routetx_req), .rrnw({\ri_rnw[1] , \ri_rnw[0] }), .a({
        \ci_a[63] , \ci_a[62] , \ci_a[61] , \ci_a[60] , \ci_a[59] , \ci_a[58] , 
        \ci_a[57] , \ci_a[56] , \ci_a[55] , \ci_a[54] , \ci_a[53] , \ci_a[52] , 
        \ci_a[51] , \ci_a[50] , \ci_a[49] , \ci_a[48] , \ci_a[47] , \ci_a[46] , 
        \ci_a[45] , \ci_a[44] , \ci_a[43] , \ci_a[42] , \ci_a[41] , \ci_a[40] , 
        \ci_a[39] , \ci_a[38] , \ci_a[37] , \ci_a[36] , \ci_a[35] , \ci_a[34] , 
        \ci_a[33] , \ci_a[32] , \ci_a[31] , \ci_a[30] , \ci_a[29] , \ci_a[28] , 
        \ci_a[27] , \ci_a[26] , \ci_a[25] , \ci_a[24] , \ci_a[23] , \ci_a[22] , 
        \ci_a[21] , \ci_a[20] , \ci_a[19] , \ci_a[18] , \ci_a[17] , \ci_a[16] , 
        \ci_a[15] , \ci_a[14] , \ci_a[13] , \ci_a[12] , \ci_a[11] , \ci_a[10] , 
        \ci_a[9] , \ci_a[8] , \ci_a[7] , \ci_a[6] , \ci_a[5] , \ci_a[4] , 
        \ci_a[3] , \ci_a[2] , \ci_a[1] , \ci_a[0] }), .chainresponse(
        chainresponse), .col({\ci_col[5] , \ci_col[4] , \ci_col[3] , 
        \ci_col[2] , \ci_col[1] , \ci_col[0] }), .crnw({\ci_rnw[1] , 
        \ci_rnw[0] }), .itag({\ci_itag[9] , \ci_itag[8] , \ci_itag[7] , 
        \ci_itag[6] , \ci_itag[5] , \ci_itag[4] , \ci_itag[3] , \ci_itag[2] , 
        \ci_itag[1] , \ci_itag[0] }), .lock({\ci_lock[1] , \ci_lock[0] }), 
        .nReset(nReset), .nchaincommandack(nchaincommandack), .pred({
        \ci_pred[1] , \ci_pred[0] }), .rack(ri_ack), .route({\route[4] , 1'b0, 
        1'b0, \route[1] , \route[0] }), .routetxack(routetx_ack), .seq({
        \ci_seq[1] , \ci_seq[0] }), .size({\ci_size[3] , \ci_size[2] , 
        \ci_size[1] , \ci_size[0] }), .wd({\ci_wd[63] , \ci_wd[62] , 
        \ci_wd[61] , \ci_wd[60] , \ci_wd[59] , \ci_wd[58] , \ci_wd[57] , 
        \ci_wd[56] , \ci_wd[55] , \ci_wd[54] , \ci_wd[53] , \ci_wd[52] , 
        \ci_wd[51] , \ci_wd[50] , \ci_wd[49] , \ci_wd[48] , \ci_wd[47] , 
        \ci_wd[46] , \ci_wd[45] , \ci_wd[44] , \ci_wd[43] , \ci_wd[42] , 
        \ci_wd[41] , \ci_wd[40] , \ci_wd[39] , \ci_wd[38] , \ci_wd[37] , 
        \ci_wd[36] , \ci_wd[35] , \ci_wd[34] , \ci_wd[33] , \ci_wd[32] , 
        \ci_wd[31] , \ci_wd[30] , \ci_wd[29] , \ci_wd[28] , \ci_wd[27] , 
        \ci_wd[26] , \ci_wd[25] , \ci_wd[24] , \ci_wd[23] , \ci_wd[22] , 
        \ci_wd[21] , \ci_wd[20] , \ci_wd[19] , \ci_wd[18] , \ci_wd[17] , 
        \ci_wd[16] , \ci_wd[15] , \ci_wd[14] , \ci_wd[13] , \ci_wd[12] , 
        \ci_wd[11] , \ci_wd[10] , \ci_wd[9] , \ci_wd[8] , \ci_wd[7] , 
        \ci_wd[6] , \ci_wd[5] , \ci_wd[4] , \ci_wd[3] , \ci_wd[2] , \ci_wd[1] , 
        \ci_wd[0] }) );
endmodule


module i_adec_tic ( e_h, e_l, r_h, r_l, ah, al, e_bare, e_dm, e_im, e_wish, 
    r_bare, r_dm, r_im, r_wish, force_bare );
output [3:0] e_h;
output [3:0] e_l;
output [3:0] r_h;
output [3:0] r_l;
input  [31:0] ah;
input  [31:0] al;
input  [3:0] e_bare;
input  [3:0] e_dm;
input  [3:0] e_im;
input  [3:0] e_wish;
input  [3:0] r_bare;
input  [3:0] r_dm;
input  [3:0] r_im;
input  [3:0] r_wish;
input  force_bare;
    wire \e_l[2] , \e_h[0] , n14, n15, \r_l[2] , \r_l[0] , im_i, dm_i, wish_i, 
        bare_i, n1, n2, n3, n6, n7, \e_l[3] , \e_l[0] , n12;
    assign e_h[3] = 1'b0;
    assign e_h[0] = \e_h[0] ;
    assign e_l[3] = \e_l[3] ;
    assign e_l[2] = \e_l[2] ;
    assign e_l[0] = \e_l[0] ;
    assign r_h[3] = \e_l[2] ;
    assign r_h[2] = \e_h[0] ;
    assign r_h[0] = 1'b0;
    assign r_l[2] = \e_l[0] ;
    assign r_l[0] = \e_l[3] ;
    ao222_1 \U1632/U18/U1/U1  ( .x(wish_i), .a(n6), .b(al[30]), .c(n6), .d(
        wish_i), .e(al[30]), .f(wish_i) );
    ao222_1 \U1633/U18/U1/U1  ( .x(bare_i), .a(n6), .b(ah[30]), .c(n6), .d(
        bare_i), .e(ah[30]), .f(bare_i) );
    ao222_1 \U1634/U18/U1/U1  ( .x(im_i), .a(al[11]), .b(n7), .c(al[11]), .d(
        im_i), .e(n7), .f(im_i) );
    ao222_1 \U1635/U18/U1/U1  ( .x(dm_i), .a(ah[11]), .b(n7), .c(ah[11]), .d(
        dm_i), .e(n7), .f(dm_i) );
    or3_1 U1 ( .x(\r_l[2] ), .a(wish_i), .b(bare_i), .c(force_bare) );
    or2_1 U2 ( .x(r_l[1]), .a(\e_l[0] ), .b(im_i) );
    or2_1 U3 ( .x(\r_l[0] ), .a(dm_i), .b(r_l[1]) );
    nor2_0 U4 ( .x(n1), .a(bare_i), .b(force_bare) );
    aoi21_1 U6 ( .x(n2), .a(n3), .b(im_i), .c(r_h[1]) );
    inv_0 U8 ( .x(n3), .a(force_bare) );
    nor2i_0 U9 ( .x(n15), .a(wish_i), .b(force_bare) );
    nor2i_0 U10 ( .x(n14), .a(dm_i), .b(force_bare) );
    inv_0 U11 ( .x(e_h[1]), .a(n1) );
    buf_1 U15 ( .x(n6), .a(ah[31]) );
    buf_1 U16 ( .x(n7), .a(al[31]) );
    nand2_2 U17 ( .x(\e_l[2] ), .a(n2), .b(n1) );
    buf_1 U18 ( .x(r_h[1]), .a(n14) );
    inv_2 U19 ( .x(\e_h[0] ), .a(n2) );
    buf_3 U20 ( .x(\e_l[3] ), .a(\r_l[0] ) );
    buf_3 U21 ( .x(\e_l[0] ), .a(\r_l[2] ) );
    nand2i_2 U22 ( .x(e_l[1]), .a(n12), .b(n2) );
    buf_1 U23 ( .x(e_h[2]), .a(n15) );
    buf_1 U24 ( .x(r_l[3]), .a(n15) );
    buf_1 U25 ( .x(n12), .a(n15) );
endmodule


module chain_selement_ga_12 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_8 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[1] , \c[0] ;
    chain_selement_ga_12 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_13 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_9 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[1] , \c[0] ;
    chain_selement_ga_13 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_14 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_10 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[1] , \c[0] ;
    chain_selement_ga_14 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_15 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_11 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[1] , \c[0] ;
    chain_selement_ga_15 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_79 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_tx_tic ( o, rtxack, e_h, e_l, noa, r_h, r_l, rtxreq );
output [4:0] o;
input  [3:0] e_h;
input  [3:0] e_l;
input  [3:0] r_h;
input  [3:0] r_l;
input  noa, rtxreq;
output rtxack;
    wire \net52[0] , \net52[1] , \net55[0] , \net55[1] , \r3[2] , \r3[1] , 
        \r3[0] , \r0[2] , \r0[1] , \r0[0] , \r2[2] , \r2[1] , \r2[0] , 
        \last[0] , \last[1] , \last[2] , \last[3] , \last[4] , \r1[2] , 
        \r1[1] , \r1[0] , net6, eopsym, net9, net11, net16, net33, net60, 
        net40, net47, net50, \I8/nb , \I8/na , \I11/nc , \I11/nb , \I11/na , 
        \I7_0_/U25/U1/clr , \I7_0_/U25/U1/ob , \I7_1_/U25/U1/clr , 
        \I7_1_/U25/U1/ob ;
    assign o[3] = 1'b0;
    assign o[2] = 1'b0;
    route_symbol_8 I0 ( .o({\r3[2] , \r3[1] , \r3[0] }), .txack(net33), 
        .txack_last(\last[4] ), .e({e_h[3], e_l[3]}), .oa(net60), .r({r_h[3], 
        r_l[3]}), .txreq(rtxreq) );
    route_symbol_9 I1 ( .o({\r2[2] , \r2[1] , \r2[0] }), .txack(net40), 
        .txack_last(\last[3] ), .e({e_h[2], e_l[2]}), .oa(net60), .r({r_h[2], 
        r_l[2]}), .txreq(net33) );
    route_symbol_10 I2 ( .o({\r1[2] , \r1[1] , \r1[0] }), .txack(net47), 
        .txack_last(\last[2] ), .e({e_h[1], e_l[1]}), .oa(net60), .r({r_h[1], 
        r_l[1]}), .txreq(net40) );
    route_symbol_11 I3 ( .o({\r0[2] , \r0[1] , \r0[0] }), .txack(net50), 
        .txack_last(\last[1] ), .e({e_h[0], e_l[0]}), .oa(net60), .r({r_h[0], 
        r_l[0]}), .txreq(net47) );
    chain_selement_ga_79 I9 ( .Aa(\last[0] ), .Br(eopsym), .Ar(net50), .Ba(
        net60) );
    nor3_1 \I8/U27  ( .x(\I8/nb ), .a(o[4]), .b(o[3]), .c(o[2]) );
    nor2_1 \I8/U26  ( .x(\I8/na ), .a(o[1]), .b(o[0]) );
    nand2_2 \I8/U29  ( .x(net60), .a(\I8/nb ), .b(\I8/na ) );
    or2_1 \I13_0_/U12  ( .x(\net55[1] ), .a(\r1[0] ), .b(\r0[0] ) );
    or2_1 \I13_1_/U12  ( .x(\net55[0] ), .a(\r1[1] ), .b(\r0[1] ) );
    or2_1 \I14_0_/U12  ( .x(\net52[1] ), .a(\r3[0] ), .b(\r2[0] ) );
    or2_1 \I14_1_/U12  ( .x(\net52[0] ), .a(\r3[1] ), .b(\r2[1] ) );
    nand3_1 \I11/U31  ( .x(rtxack), .a(\I11/nc ), .b(\I11/nb ), .c(\I11/na )
         );
    inv_1 \I11/U33  ( .x(\I11/nc ), .a(\last[0] ) );
    nor2_1 \I11/U26  ( .x(\I11/na ), .a(\last[3] ), .b(\last[4] ) );
    nor2_1 \I11/U32  ( .x(\I11/nb ), .a(\last[1] ), .b(\last[2] ) );
    nor2_1 \I16/U5  ( .x(net16), .a(\r1[2] ), .b(\r0[2] ) );
    nor2_1 \I5/U5  ( .x(net11), .a(\r3[2] ), .b(\r2[2] ) );
    nand3_1 \I17/U9  ( .x(net9), .a(net6), .b(net11), .c(net16) );
    inv_1 \I18/U3  ( .x(net6), .a(eopsym) );
    oa31_1 \I7_0_/U25/U1/Uclr  ( .x(\I7_0_/U25/U1/clr ), .a(noa), .b(
        \net55[1] ), .c(\net52[1] ), .d(o[0]) );
    oaoi211_1 \I7_0_/U25/U1/Uaoi  ( .x(\I7_0_/U25/U1/ob ), .a(\net55[1] ), .b(
        \net52[1] ), .c(noa), .d(\I7_0_/U25/U1/clr ) );
    inv_2 \I7_0_/U25/U1/Ui  ( .x(o[0]), .a(\I7_0_/U25/U1/ob ) );
    oa31_1 \I7_1_/U25/U1/Uclr  ( .x(\I7_1_/U25/U1/clr ), .a(noa), .b(
        \net55[0] ), .c(\net52[0] ), .d(o[1]) );
    oaoi211_1 \I7_1_/U25/U1/Uaoi  ( .x(\I7_1_/U25/U1/ob ), .a(\net55[0] ), .b(
        \net52[0] ), .c(noa), .d(\I7_1_/U25/U1/clr ) );
    inv_2 \I7_1_/U25/U1/Ui  ( .x(o[1]), .a(\I7_1_/U25/U1/ob ) );
    ao222_1 \I15/U18/U1/U1  ( .x(o[4]), .a(noa), .b(net9), .c(noa), .d(o[4]), 
        .e(net9), .f(o[4]) );
endmodule


module chain_dr8bit_completion_32 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_33 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_34 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_35 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr32bit_completion_6 ( o, i );
input  [63:0] i;
output o;
    wire nx, \cd[3] , \cd[2] , ny, \cd[0] , \cd[1] , \U16/Z , \U6/Z , \U15/Z ;
    chain_dr8bit_completion_32 U11 ( .o(\cd[3] ), .i({i[63], i[62], i[61], 
        i[60], i[59], i[58], i[57], i[56], i[31], i[30], i[29], i[28], i[27], 
        i[26], i[25], i[24]}) );
    chain_dr8bit_completion_35 U14 ( .o(\cd[2] ), .i({i[55], i[54], i[53], 
        i[52], i[51], i[50], i[49], i[48], i[23], i[22], i[21], i[20], i[19], 
        i[18], i[17], i[16]}) );
    chain_dr8bit_completion_34 U13 ( .o(\cd[1] ), .i({i[47], i[46], i[45], 
        i[44], i[43], i[42], i[41], i[40], i[15], i[14], i[13], i[12], i[11], 
        i[10], i[9], i[8]}) );
    chain_dr8bit_completion_33 U12 ( .o(\cd[0] ), .i({i[39], i[38], i[37], 
        i[36], i[35], i[34], i[33], i[32], i[7], i[6], i[5], i[4], i[3], i[2], 
        i[1], i[0]}) );
    aoi222_1 \U16/U30/U1  ( .x(ny), .a(\cd[0] ), .b(\cd[1] ), .c(\cd[0] ), .d(
        \U16/Z ), .e(\cd[1] ), .f(\U16/Z ) );
    inv_1 \U16/U30/Uinv  ( .x(\U16/Z ), .a(ny) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(ny), .b(nx), .c(ny), .d(\U6/Z ), .e(nx), 
        .f(\U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U15/U30/U1  ( .x(nx), .a(\cd[3] ), .b(\cd[2] ), .c(\cd[3] ), .d(
        \U15/Z ), .e(\cd[2] ), .f(\U15/Z ) );
    inv_1 \U15/U30/Uinv  ( .x(\U15/Z ), .a(nx) );
endmodule


module chain_dr8bit_completion_36 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_37 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_38 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_39 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr32bit_completion_7 ( o, i );
input  [63:0] i;
output o;
    wire nx, \cd[3] , \cd[2] , ny, \cd[0] , \cd[1] , \U16/Z , \U6/Z , \U15/Z ;
    chain_dr8bit_completion_36 U11 ( .o(\cd[3] ), .i({i[63], i[62], i[61], 
        i[60], i[59], i[58], i[57], i[56], i[31], i[30], i[29], i[28], i[27], 
        i[26], i[25], i[24]}) );
    chain_dr8bit_completion_39 U14 ( .o(\cd[2] ), .i({i[55], i[54], i[53], 
        i[52], i[51], i[50], i[49], i[48], i[23], i[22], i[21], i[20], i[19], 
        i[18], i[17], i[16]}) );
    chain_dr8bit_completion_38 U13 ( .o(\cd[1] ), .i({i[47], i[46], i[45], 
        i[44], i[43], i[42], i[41], i[40], i[15], i[14], i[13], i[12], i[11], 
        i[10], i[9], i[8]}) );
    chain_dr8bit_completion_37 U12 ( .o(\cd[0] ), .i({i[39], i[38], i[37], 
        i[36], i[35], i[34], i[33], i[32], i[7], i[6], i[5], i[4], i[3], i[2], 
        i[1], i[0]}) );
    aoi222_1 \U16/U30/U1  ( .x(ny), .a(\cd[0] ), .b(\cd[1] ), .c(\cd[0] ), .d(
        \U16/Z ), .e(\cd[1] ), .f(\U16/Z ) );
    inv_1 \U16/U30/Uinv  ( .x(\U16/Z ), .a(ny) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(ny), .b(nx), .c(ny), .d(\U6/Z ), .e(nx), 
        .f(\U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U15/U30/U1  ( .x(nx), .a(\cd[3] ), .b(\cd[2] ), .c(\cd[3] ), .d(
        \U15/Z ), .e(\cd[2] ), .f(\U15/Z ) );
    inv_1 \U15/U30/Uinv  ( .x(\U15/Z ), .a(nx) );
endmodule


module chain_dr8bit_completion_54 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_55 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_selement_ga_52 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_53 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_54 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_55 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_56 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_57 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_58 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_59 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_60 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_61 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_icmux_2 ( ack, chainh, chainl, sendack, addr, col, itag, lock, 
    nReset, nia, pred, rnw, sendreq, seq, size, wd );
output [7:0] chainh;
output [7:0] chainl;
input  [63:0] addr;
input  [5:0] col;
input  [9:0] itag;
input  [1:0] lock;
input  [1:0] pred;
input  [1:0] rnw;
input  [1:0] seq;
input  [3:0] size;
input  [63:0] wd;
input  nReset, nia, sendreq;
output ack, sendack;
    wire \net207[0] , \net207[1] , \net207[2] , \net207[3] , \net207[4] , 
        \net207[5] , \net207[6] , \net207[7] , \net207[8] , \net207[9] , 
        \net207[10] , \net207[11] , \net207[12] , \net207[13] , \net207[14] , 
        \net207[15] , \bs[0] , \bs[1] , \bs[2] , \bs[3] , \bs[4] , \bs[5] , 
        \bs[6] , \bs[7] , \bs[8] , \net231[0] , \net231[1] , \net231[2] , 
        \net231[3] , \net231[4] , \net231[5] , \net231[6] , \net231[7] , 
        \net231[8] , \net231[9] , \net231[10] , \net231[11] , \net231[12] , 
        \net231[13] , \net231[14] , \net231[15] , \hdr[4] , \net234[0] , 
        \net234[1] , \net234[2] , \net234[3] , \net234[4] , \net234[5] , 
        \net234[6] , \net234[7] , \net234[8] , \net234[9] , \net234[10] , 
        \net234[11] , \net234[12] , \net234[13] , \net234[14] , \net234[15] , 
        \net217[0] , \net217[1] , \net217[2] , \net217[3] , \net217[4] , 
        \net217[5] , \net217[6] , \net217[7] , \net217[8] , \net217[9] , 
        \net217[10] , \net217[11] , \net217[12] , \net217[13] , \net217[14] , 
        \net217[15] , \net246[0] , \net246[1] , \net246[2] , \net246[3] , 
        \net246[4] , \net246[5] , \net246[6] , \net246[7] , \net246[8] , 
        \net246[9] , \net246[10] , \net246[11] , \net246[12] , \net246[13] , 
        \net246[14] , \net246[15] , \net243[0] , \net243[1] , \net243[2] , 
        \net243[3] , \net243[4] , \net243[5] , \net243[6] , \net243[7] , 
        \net243[8] , \net243[9] , \net243[10] , \net243[11] , \net243[12] , 
        \net243[13] , \net243[14] , \net243[15] , \net240[0] , \net240[1] , 
        \net240[2] , \net240[3] , \net240[4] , \net240[5] , \net240[6] , 
        \net240[7] , \net240[8] , \net240[9] , \net240[10] , \net240[11] , 
        \net240[12] , \net240[13] , \net240[14] , \net240[15] , \net219[0] , 
        \net219[1] , \net219[2] , \net219[3] , \net219[4] , \net219[5] , 
        \net219[6] , \net219[7] , \net219[8] , \net219[9] , \net219[10] , 
        \net219[11] , \net219[12] , \net219[13] , \net219[14] , \net219[15] , 
        \net237[0] , \net237[1] , \net237[2] , \net237[5] , \net237[6] , 
        \net237[7] , \net237[8] , \net237[9] , \net237[10] , \net237[11] , 
        \net237[12] , \net237[13] , \net237[14] , \net237[15] , \net222[0] , 
        \net222[1] , \net222[2] , \net222[3] , \net222[4] , \net222[5] , 
        \net222[6] , \net222[7] , \net222[8] , \net222[9] , \net222[10] , 
        \net222[11] , \net222[12] , \net222[13] , \net222[14] , \net222[15] , 
        \net225[0] , \net225[1] , \net225[2] , \net225[3] , \net225[4] , 
        \net225[5] , \net225[6] , \net225[7] , \net225[8] , \net225[9] , 
        \net225[10] , \net225[11] , \net225[12] , \net225[13] , \net225[14] , 
        \net225[15] , \net228[0] , \net228[1] , \net228[2] , \net228[3] , 
        \net228[4] , \net228[5] , \net228[6] , \net228[7] , \net228[8] , 
        \net228[9] , \net228[10] , \net228[11] , \net228[12] , \net228[13] , 
        \net228[14] , \net228[15] , \net212[0] , \net212[1] , \net212[2] , 
        \net212[3] , \net212[4] , \net212[5] , \net212[6] , \net212[7] , 
        \net212[8] , \net212[9] , \net212[10] , \net212[11] , \net212[12] , 
        \net212[13] , \net212[14] , \net212[15] , net138, net198, net176, 
        net132, net131, net136, net185, net187, net191, net293, net152, net146, 
        net148, net156, net160, net168, net172, net164, net289, net180, net189, 
        net249, net261, net251, net255, net253, net259, net269, net267, net263, 
        net265, \U40_0_/n5 , \U40_0_/n3 , \U40_0_/n4 , \U40_1_/n5 , 
        \U40_1_/n3 , \U40_1_/n4 , \U40_2_/n5 , \U40_2_/n3 , \U40_2_/n4 , 
        \U40_3_/n5 , \U40_3_/n3 , \U40_3_/n4 , \U40_4_/n5 , \U40_4_/n3 , 
        \U40_4_/n4 , \U40_5_/n5 , \U40_5_/n3 , \U40_5_/n4 , \U40_6_/n5 , 
        \U40_6_/n3 , \U40_6_/n4 , \U40_7_/n5 , \U40_7_/n3 , \U40_7_/n4 , 
        \U40_8_/n5 , \U40_8_/n3 , \U40_8_/n4 , \U40_9_/n5 , \U40_9_/n3 , 
        \U40_9_/n4 , \U40_10_/n5 , \U40_10_/n3 , \U40_10_/n4 , \U40_11_/n5 , 
        \U40_11_/n3 , \U40_11_/n4 , \U40_12_/n5 , \U40_12_/n3 , \U40_12_/n4 , 
        \U40_13_/n5 , \U40_13_/n3 , \U40_13_/n4 , \U40_14_/n5 , \U40_14_/n3 , 
        \U40_14_/n4 , \U40_15_/n5 , \U40_15_/n3 , \U40_15_/n4 , \U14_0_/n5 , 
        \U14_0_/n1 , \U14_0_/n2 , \U14_0_/n3 , \U14_0_/n4 , \U14_1_/n5 , 
        \U14_1_/n1 , \U14_1_/n2 , \U14_1_/n3 , \U14_1_/n4 , \U14_2_/n5 , 
        \U14_2_/n1 , \U14_2_/n2 , \U14_2_/n3 , \U14_2_/n4 , \U14_3_/n5 , 
        \U14_3_/n1 , \U14_3_/n2 , \U14_3_/n3 , \U14_3_/n4 , \U14_4_/n5 , 
        \U14_4_/n1 , \U14_4_/n2 , \U14_4_/n3 , \U14_4_/n4 , \U14_5_/n5 , 
        \U14_5_/n1 , \U14_5_/n2 , \U14_5_/n3 , \U14_5_/n4 , \U14_6_/n5 , 
        \U14_6_/n1 , \U14_6_/n2 , \U14_6_/n3 , \U14_6_/n4 , \U14_7_/n5 , 
        \U14_7_/n1 , \U14_7_/n2 , \U14_7_/n3 , \U14_7_/n4 , \U14_8_/n5 , 
        \U14_8_/n1 , \U14_8_/n2 , \U14_8_/n3 , \U14_8_/n4 , \U14_9_/n5 , 
        \U14_9_/n1 , \U14_9_/n2 , \U14_9_/n3 , \U14_9_/n4 , \U14_10_/n5 , 
        \U14_10_/n1 , \U14_10_/n2 , \U14_10_/n3 , \U14_10_/n4 , \U14_11_/n5 , 
        \U14_11_/n1 , \U14_11_/n2 , \U14_11_/n4 , \U14_12_/n5 , \U14_12_/n1 , 
        \U14_12_/n2 , \U14_12_/n4 , \U14_13_/n5 , \U14_13_/n1 , \U14_13_/n2 , 
        \U14_13_/n3 , \U14_13_/n4 , \U14_14_/n5 , \U14_14_/n1 , \U14_14_/n2 , 
        \U14_14_/n3 , \U14_14_/n4 , \U14_15_/n5 , \U14_15_/n1 , \U14_15_/n2 , 
        \U14_15_/n3 , \U14_15_/n4 , \U91_0_/n5 , \U91_0_/n1 , \U91_0_/n2 , 
        \U91_0_/n3 , \U91_0_/n4 , \U91_1_/n5 , \U91_1_/n1 , \U91_1_/n2 , 
        \U91_1_/n3 , \U91_1_/n4 , \U91_2_/n5 , \U91_2_/n1 , \U91_2_/n2 , 
        \U91_2_/n3 , \U91_2_/n4 , \U91_3_/n5 , \U91_3_/n1 , \U91_3_/n2 , 
        \U91_3_/n3 , \U91_3_/n4 , \U91_4_/n5 , \U91_4_/n1 , \U91_4_/n2 , 
        \U91_4_/n3 , \U91_4_/n4 , \U91_5_/n5 , \U91_5_/n1 , \U91_5_/n2 , 
        \U91_5_/n3 , \U91_5_/n4 , \U91_6_/n5 , \U91_6_/n1 , \U91_6_/n2 , 
        \U91_6_/n3 , \U91_6_/n4 , \U91_7_/n5 , \U91_7_/n1 , \U91_7_/n2 , 
        \U91_7_/n3 , \U91_7_/n4 , \U91_8_/n5 , \U91_8_/n1 , \U91_8_/n2 , 
        \U91_8_/n3 , \U91_8_/n4 , \U91_9_/n5 , \U91_9_/n1 , \U91_9_/n2 , 
        \U91_9_/n3 , \U91_9_/n4 , \U91_10_/n5 , \U91_10_/n1 , \U91_10_/n2 , 
        \U91_10_/n3 , \U91_10_/n4 , \U91_11_/n5 , \U91_11_/n1 , \U91_11_/n2 , 
        \U91_11_/n3 , \U91_11_/n4 , \U91_12_/n5 , \U91_12_/n1 , \U91_12_/n2 , 
        \U91_12_/n3 , \U91_12_/n4 , \U91_13_/n5 , \U91_13_/n1 , \U91_13_/n2 , 
        \U91_13_/n3 , \U91_13_/n4 , \U91_14_/n5 , \U91_14_/n1 , \U91_14_/n2 , 
        \U91_14_/n3 , \U91_14_/n4 , \U91_15_/n5 , \U91_15_/n1 , \U91_15_/n2 , 
        \U91_15_/n3 , \U91_15_/n4 , \U148/U21/nr , \U148/U21/nd , 
        \U148/U21/n2 , \U151/Z , n1;
    chain_selement_ga_53 U163 ( .Aa(net152), .Br(net146), .Ar(net148), .Ba(n1)
         );
    chain_selement_ga_54 U164 ( .Aa(net156), .Br(\bs[1] ), .Ar(net152), .Ba(
        net138) );
    chain_selement_ga_55 U165 ( .Aa(net160), .Br(\bs[2] ), .Ar(net156), .Ba(n1
        ) );
    chain_selement_ga_56 U166 ( .Aa(net168), .Br(\bs[3] ), .Ar(net160), .Ba(
        net138) );
    chain_selement_ga_60 U170 ( .Aa(net172), .Br(\bs[7] ), .Ar(net164), .Ba(
        net138) );
    chain_selement_ga_57 U167 ( .Aa(net132), .Br(\bs[4] ), .Ar(net168), .Ba(
        net138) );
    chain_selement_ga_61 U171 ( .Aa(net289), .Br(\bs[8] ), .Ar(net172), .Ba(
        net138) );
    chain_selement_ga_58 U168 ( .Aa(net180), .Br(\bs[5] ), .Ar(net176), .Ba(
        net138) );
    chain_selement_ga_59 U169 ( .Aa(net164), .Br(\bs[6] ), .Ar(net180), .Ba(n1
        ) );
    chain_selement_ga_52 U161 ( .Aa(net148), .Br(\bs[0] ), .Ar(\hdr[4] ), .Ba(
        n1) );
    chain_dr8bit_completion_54 U119 ( .o(net185), .i({col[5], col[4], col[3], 
        itag[9], itag[8], itag[7], itag[6], itag[5], col[2], col[1], col[0], 
        itag[4], itag[3], itag[2], itag[1], itag[0]}) );
    chain_dr8bit_completion_55 U147 ( .o(net187), .i({size[3], size[2], rnw[1], 
        1'b0, 1'b0, lock[1], pred[1], seq[1], size[1], size[0], rnw[0], 
        \hdr[4] , \hdr[4] , lock[0], pred[0], seq[0]}) );
    chain_dr32bit_completion_6 U117 ( .o(net189), .i(wd) );
    chain_dr32bit_completion_7 U118 ( .o(net191), .i(addr) );
    or2_4 \U122/U12  ( .x(net293), .a(net189), .b(net131) );
    or2_4 \U53/U12  ( .x(sendack), .a(net131), .b(net289) );
    and2_1 \U32_0_/U8  ( .x(\net246[15] ), .a(itag[0]), .b(net265) );
    and2_1 \U32_1_/U8  ( .x(\net246[14] ), .a(itag[1]), .b(net265) );
    and2_1 \U32_2_/U8  ( .x(\net246[13] ), .a(itag[2]), .b(net265) );
    and2_1 \U32_3_/U8  ( .x(\net246[12] ), .a(itag[3]), .b(net265) );
    and2_1 \U32_4_/U8  ( .x(\net246[11] ), .a(itag[4]), .b(net265) );
    and2_1 \U32_5_/U8  ( .x(\net246[10] ), .a(col[0]), .b(net265) );
    and2_1 \U32_6_/U8  ( .x(\net246[9] ), .a(col[1]), .b(net265) );
    and2_1 \U32_7_/U8  ( .x(\net246[8] ), .a(col[2]), .b(net265) );
    and2_1 \U32_8_/U8  ( .x(\net246[7] ), .a(itag[5]), .b(net265) );
    and2_1 \U32_9_/U8  ( .x(\net246[6] ), .a(itag[6]), .b(net265) );
    and2_1 \U32_10_/U8  ( .x(\net246[5] ), .a(itag[7]), .b(net265) );
    and2_1 \U32_11_/U8  ( .x(\net246[4] ), .a(itag[8]), .b(net265) );
    and2_1 \U32_12_/U8  ( .x(\net246[3] ), .a(itag[9]), .b(net265) );
    and2_1 \U32_13_/U8  ( .x(\net246[2] ), .a(col[3]), .b(net265) );
    and2_1 \U32_14_/U8  ( .x(\net246[1] ), .a(col[4]), .b(net265) );
    and2_1 \U32_15_/U8  ( .x(\net246[0] ), .a(col[5]), .b(net265) );
    and2_1 \U76_0_/U8  ( .x(\net243[15] ), .a(wd[8]), .b(net263) );
    and2_1 \U76_1_/U8  ( .x(\net243[14] ), .a(wd[9]), .b(net263) );
    and2_1 \U76_2_/U8  ( .x(\net243[13] ), .a(wd[10]), .b(net263) );
    and2_1 \U76_3_/U8  ( .x(\net243[12] ), .a(wd[11]), .b(net263) );
    and2_1 \U76_4_/U8  ( .x(\net243[11] ), .a(wd[12]), .b(net263) );
    and2_1 \U76_5_/U8  ( .x(\net243[10] ), .a(wd[13]), .b(net263) );
    and2_1 \U76_6_/U8  ( .x(\net243[9] ), .a(wd[14]), .b(net263) );
    and2_1 \U76_7_/U8  ( .x(\net243[8] ), .a(wd[15]), .b(net263) );
    and2_1 \U76_8_/U8  ( .x(\net243[7] ), .a(wd[40]), .b(net263) );
    and2_1 \U76_9_/U8  ( .x(\net243[6] ), .a(wd[41]), .b(net263) );
    and2_1 \U76_10_/U8  ( .x(\net243[5] ), .a(wd[42]), .b(net263) );
    and2_1 \U76_11_/U8  ( .x(\net243[4] ), .a(wd[43]), .b(net263) );
    and2_1 \U76_12_/U8  ( .x(\net243[3] ), .a(wd[44]), .b(net263) );
    and2_1 \U76_13_/U8  ( .x(\net243[2] ), .a(wd[45]), .b(net263) );
    and2_1 \U76_14_/U8  ( .x(\net243[1] ), .a(wd[46]), .b(net263) );
    and2_1 \U76_15_/U8  ( .x(\net243[0] ), .a(wd[47]), .b(net263) );
    and2_1 \U80_0_/U8  ( .x(\net240[15] ), .a(wd[16]), .b(net267) );
    and2_1 \U80_1_/U8  ( .x(\net240[14] ), .a(wd[17]), .b(net267) );
    and2_1 \U80_2_/U8  ( .x(\net240[13] ), .a(wd[18]), .b(net267) );
    and2_1 \U80_3_/U8  ( .x(\net240[12] ), .a(wd[19]), .b(net267) );
    and2_1 \U80_4_/U8  ( .x(\net240[11] ), .a(wd[20]), .b(net267) );
    and2_1 \U80_5_/U8  ( .x(\net240[10] ), .a(wd[21]), .b(net267) );
    and2_1 \U80_6_/U8  ( .x(\net240[9] ), .a(wd[22]), .b(net267) );
    and2_1 \U80_7_/U8  ( .x(\net240[8] ), .a(wd[23]), .b(net267) );
    and2_1 \U80_8_/U8  ( .x(\net240[7] ), .a(wd[48]), .b(net267) );
    and2_1 \U80_9_/U8  ( .x(\net240[6] ), .a(wd[49]), .b(net267) );
    and2_1 \U80_10_/U8  ( .x(\net240[5] ), .a(wd[50]), .b(net267) );
    and2_1 \U80_11_/U8  ( .x(\net240[4] ), .a(wd[51]), .b(net267) );
    and2_1 \U80_12_/U8  ( .x(\net240[3] ), .a(wd[52]), .b(net267) );
    and2_1 \U80_13_/U8  ( .x(\net240[2] ), .a(wd[53]), .b(net267) );
    and2_1 \U80_14_/U8  ( .x(\net240[1] ), .a(wd[54]), .b(net267) );
    and2_1 \U80_15_/U8  ( .x(\net240[0] ), .a(wd[55]), .b(net267) );
    and2_1 \U128_0_/U8  ( .x(\net237[15] ), .a(seq[0]), .b(net269) );
    and2_1 \U128_1_/U8  ( .x(\net237[14] ), .a(pred[0]), .b(net269) );
    and2_1 \U128_2_/U8  ( .x(\net237[13] ), .a(lock[0]), .b(net269) );
    and2_1 \U128_3_/U8  ( .x(\net237[12] ), .a(\hdr[4] ), .b(net269) );
    and2_1 \U128_4_/U8  ( .x(\net237[11] ), .a(\hdr[4] ), .b(net269) );
    and2_1 \U128_5_/U8  ( .x(\net237[10] ), .a(rnw[0]), .b(net269) );
    and2_1 \U128_6_/U8  ( .x(\net237[9] ), .a(size[0]), .b(net269) );
    and2_1 \U128_7_/U8  ( .x(\net237[8] ), .a(size[1]), .b(net269) );
    and2_1 \U128_8_/U8  ( .x(\net237[7] ), .a(seq[1]), .b(net269) );
    and2_1 \U128_9_/U8  ( .x(\net237[6] ), .a(pred[1]), .b(net269) );
    and2_1 \U128_10_/U8  ( .x(\net237[5] ), .a(lock[1]), .b(net269) );
    and2_1 \U128_13_/U8  ( .x(\net237[2] ), .a(rnw[1]), .b(net269) );
    and2_1 \U128_14_/U8  ( .x(\net237[1] ), .a(size[2]), .b(net269) );
    and2_1 \U128_15_/U8  ( .x(\net237[0] ), .a(size[3]), .b(net269) );
    and2_1 \U37_0_/U8  ( .x(\net234[15] ), .a(addr[8]), .b(net259) );
    and2_1 \U37_1_/U8  ( .x(\net234[14] ), .a(addr[9]), .b(net259) );
    and2_1 \U37_2_/U8  ( .x(\net234[13] ), .a(addr[10]), .b(net259) );
    and2_1 \U37_3_/U8  ( .x(\net234[12] ), .a(addr[11]), .b(net259) );
    and2_1 \U37_4_/U8  ( .x(\net234[11] ), .a(addr[12]), .b(net259) );
    and2_1 \U37_5_/U8  ( .x(\net234[10] ), .a(addr[13]), .b(net259) );
    and2_1 \U37_6_/U8  ( .x(\net234[9] ), .a(addr[14]), .b(net259) );
    and2_1 \U37_7_/U8  ( .x(\net234[8] ), .a(addr[15]), .b(net259) );
    and2_1 \U37_8_/U8  ( .x(\net234[7] ), .a(addr[40]), .b(net259) );
    and2_1 \U37_9_/U8  ( .x(\net234[6] ), .a(addr[41]), .b(net259) );
    and2_1 \U37_10_/U8  ( .x(\net234[5] ), .a(addr[42]), .b(net259) );
    and2_1 \U37_11_/U8  ( .x(\net234[4] ), .a(addr[43]), .b(net259) );
    and2_1 \U37_12_/U8  ( .x(\net234[3] ), .a(addr[44]), .b(net259) );
    and2_1 \U37_13_/U8  ( .x(\net234[2] ), .a(addr[45]), .b(net259) );
    and2_1 \U37_14_/U8  ( .x(\net234[1] ), .a(addr[46]), .b(net259) );
    and2_1 \U37_15_/U8  ( .x(\net234[0] ), .a(addr[47]), .b(net259) );
    and2_1 \U33_0_/U8  ( .x(\net231[15] ), .a(addr[16]), .b(net253) );
    and2_1 \U33_1_/U8  ( .x(\net231[14] ), .a(addr[17]), .b(net253) );
    and2_1 \U33_2_/U8  ( .x(\net231[13] ), .a(addr[18]), .b(net253) );
    and2_1 \U33_3_/U8  ( .x(\net231[12] ), .a(addr[19]), .b(net253) );
    and2_1 \U33_4_/U8  ( .x(\net231[11] ), .a(addr[20]), .b(net253) );
    and2_1 \U33_5_/U8  ( .x(\net231[10] ), .a(addr[21]), .b(net253) );
    and2_1 \U33_6_/U8  ( .x(\net231[9] ), .a(addr[22]), .b(net253) );
    and2_1 \U33_7_/U8  ( .x(\net231[8] ), .a(addr[23]), .b(net253) );
    and2_1 \U33_8_/U8  ( .x(\net231[7] ), .a(addr[48]), .b(net253) );
    and2_1 \U33_9_/U8  ( .x(\net231[6] ), .a(addr[49]), .b(net253) );
    and2_1 \U33_10_/U8  ( .x(\net231[5] ), .a(addr[50]), .b(net253) );
    and2_1 \U33_11_/U8  ( .x(\net231[4] ), .a(addr[51]), .b(net253) );
    and2_1 \U33_12_/U8  ( .x(\net231[3] ), .a(addr[52]), .b(net253) );
    and2_1 \U33_13_/U8  ( .x(\net231[2] ), .a(addr[53]), .b(net253) );
    and2_1 \U33_14_/U8  ( .x(\net231[1] ), .a(addr[54]), .b(net253) );
    and2_1 \U33_15_/U8  ( .x(\net231[0] ), .a(addr[55]), .b(net253) );
    and2_1 \U81_0_/U8  ( .x(\net228[15] ), .a(wd[24]), .b(net255) );
    and2_1 \U81_1_/U8  ( .x(\net228[14] ), .a(wd[25]), .b(net255) );
    and2_1 \U81_2_/U8  ( .x(\net228[13] ), .a(wd[26]), .b(net255) );
    and2_1 \U81_3_/U8  ( .x(\net228[12] ), .a(wd[27]), .b(net255) );
    and2_1 \U81_4_/U8  ( .x(\net228[11] ), .a(wd[28]), .b(net255) );
    and2_1 \U81_5_/U8  ( .x(\net228[10] ), .a(wd[29]), .b(net255) );
    and2_1 \U81_6_/U8  ( .x(\net228[9] ), .a(wd[30]), .b(net255) );
    and2_1 \U81_7_/U8  ( .x(\net228[8] ), .a(wd[31]), .b(net255) );
    and2_1 \U81_8_/U8  ( .x(\net228[7] ), .a(wd[56]), .b(net255) );
    and2_1 \U81_9_/U8  ( .x(\net228[6] ), .a(wd[57]), .b(net255) );
    and2_1 \U81_10_/U8  ( .x(\net228[5] ), .a(wd[58]), .b(net255) );
    and2_1 \U81_11_/U8  ( .x(\net228[4] ), .a(wd[59]), .b(net255) );
    and2_1 \U81_12_/U8  ( .x(\net228[3] ), .a(wd[60]), .b(net255) );
    and2_1 \U81_13_/U8  ( .x(\net228[2] ), .a(wd[61]), .b(net255) );
    and2_1 \U81_14_/U8  ( .x(\net228[1] ), .a(wd[62]), .b(net255) );
    and2_1 \U81_15_/U8  ( .x(\net228[0] ), .a(wd[63]), .b(net255) );
    and2_1 \U34_0_/U8  ( .x(\net225[15] ), .a(addr[0]), .b(net251) );
    and2_1 \U34_1_/U8  ( .x(\net225[14] ), .a(addr[1]), .b(net251) );
    and2_1 \U34_2_/U8  ( .x(\net225[13] ), .a(addr[2]), .b(net251) );
    and2_1 \U34_3_/U8  ( .x(\net225[12] ), .a(addr[3]), .b(net251) );
    and2_1 \U34_4_/U8  ( .x(\net225[11] ), .a(addr[4]), .b(net251) );
    and2_1 \U34_5_/U8  ( .x(\net225[10] ), .a(addr[5]), .b(net251) );
    and2_1 \U34_6_/U8  ( .x(\net225[9] ), .a(addr[6]), .b(net251) );
    and2_1 \U34_7_/U8  ( .x(\net225[8] ), .a(addr[7]), .b(net251) );
    and2_1 \U34_8_/U8  ( .x(\net225[7] ), .a(addr[32]), .b(net251) );
    and2_1 \U34_9_/U8  ( .x(\net225[6] ), .a(addr[33]), .b(net251) );
    and2_1 \U34_10_/U8  ( .x(\net225[5] ), .a(addr[34]), .b(net251) );
    and2_1 \U34_11_/U8  ( .x(\net225[4] ), .a(addr[35]), .b(net251) );
    and2_1 \U34_12_/U8  ( .x(\net225[3] ), .a(addr[36]), .b(net251) );
    and2_1 \U34_13_/U8  ( .x(\net225[2] ), .a(addr[37]), .b(net251) );
    and2_1 \U34_14_/U8  ( .x(\net225[1] ), .a(addr[38]), .b(net251) );
    and2_1 \U34_15_/U8  ( .x(\net225[0] ), .a(addr[39]), .b(net251) );
    and2_1 \U30_0_/U8  ( .x(\net222[15] ), .a(addr[24]), .b(net261) );
    and2_1 \U30_1_/U8  ( .x(\net222[14] ), .a(addr[25]), .b(net261) );
    and2_1 \U30_2_/U8  ( .x(\net222[13] ), .a(addr[26]), .b(net261) );
    and2_1 \U30_3_/U8  ( .x(\net222[12] ), .a(addr[27]), .b(net261) );
    and2_1 \U30_4_/U8  ( .x(\net222[11] ), .a(addr[28]), .b(net261) );
    and2_1 \U30_5_/U8  ( .x(\net222[10] ), .a(addr[29]), .b(net261) );
    and2_1 \U30_6_/U8  ( .x(\net222[9] ), .a(addr[30]), .b(net261) );
    and2_1 \U30_7_/U8  ( .x(\net222[8] ), .a(addr[31]), .b(net261) );
    and2_1 \U30_8_/U8  ( .x(\net222[7] ), .a(addr[56]), .b(net261) );
    and2_1 \U30_9_/U8  ( .x(\net222[6] ), .a(addr[57]), .b(net261) );
    and2_1 \U30_10_/U8  ( .x(\net222[5] ), .a(addr[58]), .b(net261) );
    and2_1 \U30_11_/U8  ( .x(\net222[4] ), .a(addr[59]), .b(net261) );
    and2_1 \U30_12_/U8  ( .x(\net222[3] ), .a(addr[60]), .b(net261) );
    and2_1 \U30_13_/U8  ( .x(\net222[2] ), .a(addr[61]), .b(net261) );
    and2_1 \U30_14_/U8  ( .x(\net222[1] ), .a(addr[62]), .b(net261) );
    and2_1 \U30_15_/U8  ( .x(\net222[0] ), .a(addr[63]), .b(net261) );
    and2_1 \U82_0_/U8  ( .x(\net219[15] ), .a(wd[0]), .b(net249) );
    and2_1 \U82_1_/U8  ( .x(\net219[14] ), .a(wd[1]), .b(net249) );
    and2_1 \U82_2_/U8  ( .x(\net219[13] ), .a(wd[2]), .b(net249) );
    and2_1 \U82_3_/U8  ( .x(\net219[12] ), .a(wd[3]), .b(net249) );
    and2_1 \U82_4_/U8  ( .x(\net219[11] ), .a(wd[4]), .b(net249) );
    and2_1 \U82_5_/U8  ( .x(\net219[10] ), .a(wd[5]), .b(net249) );
    and2_1 \U82_6_/U8  ( .x(\net219[9] ), .a(wd[6]), .b(net249) );
    and2_1 \U82_7_/U8  ( .x(\net219[8] ), .a(wd[7]), .b(net249) );
    and2_1 \U82_8_/U8  ( .x(\net219[7] ), .a(wd[32]), .b(net249) );
    and2_1 \U82_9_/U8  ( .x(\net219[6] ), .a(wd[33]), .b(net249) );
    and2_1 \U82_10_/U8  ( .x(\net219[5] ), .a(wd[34]), .b(net249) );
    and2_1 \U82_11_/U8  ( .x(\net219[4] ), .a(wd[35]), .b(net249) );
    and2_1 \U82_12_/U8  ( .x(\net219[3] ), .a(wd[36]), .b(net249) );
    and2_1 \U82_13_/U8  ( .x(\net219[2] ), .a(wd[37]), .b(net249) );
    and2_1 \U82_14_/U8  ( .x(\net219[1] ), .a(wd[38]), .b(net249) );
    and2_1 \U82_15_/U8  ( .x(\net219[0] ), .a(wd[39]), .b(net249) );
    inv_1 \U40_0_/U3  ( .x(\U40_0_/n3 ), .a(\net225[15] ) );
    inv_1 \U40_0_/U4  ( .x(\U40_0_/n4 ), .a(\net234[15] ) );
    inv_1 \U40_0_/U5  ( .x(\net217[15] ), .a(\U40_0_/n5 ) );
    inv_1 \U40_1_/U3  ( .x(\U40_1_/n3 ), .a(\net225[14] ) );
    inv_1 \U40_1_/U4  ( .x(\U40_1_/n4 ), .a(\net234[14] ) );
    inv_1 \U40_1_/U5  ( .x(\net217[14] ), .a(\U40_1_/n5 ) );
    inv_1 \U40_2_/U3  ( .x(\U40_2_/n3 ), .a(\net225[13] ) );
    inv_1 \U40_2_/U4  ( .x(\U40_2_/n4 ), .a(\net234[13] ) );
    inv_1 \U40_2_/U5  ( .x(\net217[13] ), .a(\U40_2_/n5 ) );
    inv_1 \U40_3_/U3  ( .x(\U40_3_/n3 ), .a(\net225[12] ) );
    inv_1 \U40_3_/U4  ( .x(\U40_3_/n4 ), .a(\net234[12] ) );
    inv_1 \U40_3_/U5  ( .x(\net217[12] ), .a(\U40_3_/n5 ) );
    inv_1 \U40_4_/U3  ( .x(\U40_4_/n3 ), .a(\net225[11] ) );
    inv_1 \U40_4_/U4  ( .x(\U40_4_/n4 ), .a(\net234[11] ) );
    inv_1 \U40_4_/U5  ( .x(\net217[11] ), .a(\U40_4_/n5 ) );
    inv_1 \U40_5_/U3  ( .x(\U40_5_/n3 ), .a(\net225[10] ) );
    inv_1 \U40_5_/U4  ( .x(\U40_5_/n4 ), .a(\net234[10] ) );
    inv_1 \U40_5_/U5  ( .x(\net217[10] ), .a(\U40_5_/n5 ) );
    inv_1 \U40_6_/U3  ( .x(\U40_6_/n3 ), .a(\net225[9] ) );
    inv_1 \U40_6_/U4  ( .x(\U40_6_/n4 ), .a(\net234[9] ) );
    inv_1 \U40_6_/U5  ( .x(\net217[9] ), .a(\U40_6_/n5 ) );
    inv_1 \U40_7_/U3  ( .x(\U40_7_/n3 ), .a(\net225[8] ) );
    inv_1 \U40_7_/U4  ( .x(\U40_7_/n4 ), .a(\net234[8] ) );
    inv_1 \U40_7_/U5  ( .x(\net217[8] ), .a(\U40_7_/n5 ) );
    inv_1 \U40_8_/U3  ( .x(\U40_8_/n3 ), .a(\net225[7] ) );
    inv_1 \U40_8_/U4  ( .x(\U40_8_/n4 ), .a(\net234[7] ) );
    inv_1 \U40_8_/U5  ( .x(\net217[7] ), .a(\U40_8_/n5 ) );
    inv_1 \U40_9_/U3  ( .x(\U40_9_/n3 ), .a(\net225[6] ) );
    inv_1 \U40_9_/U4  ( .x(\U40_9_/n4 ), .a(\net234[6] ) );
    inv_1 \U40_9_/U5  ( .x(\net217[6] ), .a(\U40_9_/n5 ) );
    inv_1 \U40_10_/U3  ( .x(\U40_10_/n3 ), .a(\net225[5] ) );
    inv_1 \U40_10_/U4  ( .x(\U40_10_/n4 ), .a(\net234[5] ) );
    inv_1 \U40_10_/U5  ( .x(\net217[5] ), .a(\U40_10_/n5 ) );
    inv_1 \U40_11_/U3  ( .x(\U40_11_/n3 ), .a(\net225[4] ) );
    inv_1 \U40_11_/U4  ( .x(\U40_11_/n4 ), .a(\net234[4] ) );
    inv_1 \U40_11_/U5  ( .x(\net217[4] ), .a(\U40_11_/n5 ) );
    inv_1 \U40_12_/U3  ( .x(\U40_12_/n3 ), .a(\net225[3] ) );
    inv_1 \U40_12_/U4  ( .x(\U40_12_/n4 ), .a(\net234[3] ) );
    inv_1 \U40_12_/U5  ( .x(\net217[3] ), .a(\U40_12_/n5 ) );
    inv_1 \U40_13_/U3  ( .x(\U40_13_/n3 ), .a(\net225[2] ) );
    inv_1 \U40_13_/U4  ( .x(\U40_13_/n4 ), .a(\net234[2] ) );
    inv_1 \U40_13_/U5  ( .x(\net217[2] ), .a(\U40_13_/n5 ) );
    inv_1 \U40_14_/U3  ( .x(\U40_14_/n3 ), .a(\net225[1] ) );
    inv_1 \U40_14_/U4  ( .x(\U40_14_/n4 ), .a(\net234[1] ) );
    inv_1 \U40_14_/U5  ( .x(\net217[1] ), .a(\U40_14_/n5 ) );
    inv_1 \U40_15_/U3  ( .x(\U40_15_/n3 ), .a(\net225[0] ) );
    inv_1 \U40_15_/U4  ( .x(\U40_15_/n4 ), .a(\net234[0] ) );
    inv_1 \U40_15_/U5  ( .x(\net217[0] ), .a(\U40_15_/n5 ) );
    and4_1 \U14_0_/U16  ( .x(\U14_0_/n5 ), .a(\U14_0_/n1 ), .b(\U14_0_/n2 ), 
        .c(\U14_0_/n3 ), .d(\U14_0_/n4 ) );
    inv_1 \U14_0_/U1  ( .x(\U14_0_/n1 ), .a(\net231[15] ) );
    inv_1 \U14_0_/U2  ( .x(\U14_0_/n2 ), .a(\net222[15] ) );
    inv_1 \U14_0_/U3  ( .x(\U14_0_/n3 ), .a(\net237[15] ) );
    inv_1 \U14_0_/U4  ( .x(\U14_0_/n4 ), .a(\net246[15] ) );
    inv_1 \U14_0_/U5  ( .x(\net212[15] ), .a(\U14_0_/n5 ) );
    and4_1 \U14_1_/U16  ( .x(\U14_1_/n5 ), .a(\U14_1_/n1 ), .b(\U14_1_/n2 ), 
        .c(\U14_1_/n3 ), .d(\U14_1_/n4 ) );
    inv_1 \U14_1_/U1  ( .x(\U14_1_/n1 ), .a(\net231[14] ) );
    inv_1 \U14_1_/U2  ( .x(\U14_1_/n2 ), .a(\net222[14] ) );
    inv_1 \U14_1_/U3  ( .x(\U14_1_/n3 ), .a(\net237[14] ) );
    inv_1 \U14_1_/U4  ( .x(\U14_1_/n4 ), .a(\net246[14] ) );
    inv_1 \U14_1_/U5  ( .x(\net212[14] ), .a(\U14_1_/n5 ) );
    and4_1 \U14_2_/U16  ( .x(\U14_2_/n5 ), .a(\U14_2_/n1 ), .b(\U14_2_/n2 ), 
        .c(\U14_2_/n3 ), .d(\U14_2_/n4 ) );
    inv_1 \U14_2_/U1  ( .x(\U14_2_/n1 ), .a(\net231[13] ) );
    inv_1 \U14_2_/U2  ( .x(\U14_2_/n2 ), .a(\net222[13] ) );
    inv_1 \U14_2_/U3  ( .x(\U14_2_/n3 ), .a(\net237[13] ) );
    inv_1 \U14_2_/U4  ( .x(\U14_2_/n4 ), .a(\net246[13] ) );
    inv_1 \U14_2_/U5  ( .x(\net212[13] ), .a(\U14_2_/n5 ) );
    and4_1 \U14_3_/U16  ( .x(\U14_3_/n5 ), .a(\U14_3_/n1 ), .b(\U14_3_/n2 ), 
        .c(\U14_3_/n3 ), .d(\U14_3_/n4 ) );
    inv_1 \U14_3_/U1  ( .x(\U14_3_/n1 ), .a(\net231[12] ) );
    inv_1 \U14_3_/U2  ( .x(\U14_3_/n2 ), .a(\net222[12] ) );
    inv_1 \U14_3_/U3  ( .x(\U14_3_/n3 ), .a(\net237[12] ) );
    inv_1 \U14_3_/U4  ( .x(\U14_3_/n4 ), .a(\net246[12] ) );
    inv_1 \U14_3_/U5  ( .x(\net212[12] ), .a(\U14_3_/n5 ) );
    and4_1 \U14_4_/U16  ( .x(\U14_4_/n5 ), .a(\U14_4_/n1 ), .b(\U14_4_/n2 ), 
        .c(\U14_4_/n3 ), .d(\U14_4_/n4 ) );
    inv_1 \U14_4_/U1  ( .x(\U14_4_/n1 ), .a(\net231[11] ) );
    inv_1 \U14_4_/U2  ( .x(\U14_4_/n2 ), .a(\net222[11] ) );
    inv_1 \U14_4_/U3  ( .x(\U14_4_/n3 ), .a(\net237[11] ) );
    inv_1 \U14_4_/U4  ( .x(\U14_4_/n4 ), .a(\net246[11] ) );
    inv_1 \U14_4_/U5  ( .x(\net212[11] ), .a(\U14_4_/n5 ) );
    and4_1 \U14_5_/U16  ( .x(\U14_5_/n5 ), .a(\U14_5_/n1 ), .b(\U14_5_/n2 ), 
        .c(\U14_5_/n3 ), .d(\U14_5_/n4 ) );
    inv_1 \U14_5_/U1  ( .x(\U14_5_/n1 ), .a(\net231[10] ) );
    inv_1 \U14_5_/U2  ( .x(\U14_5_/n2 ), .a(\net222[10] ) );
    inv_1 \U14_5_/U3  ( .x(\U14_5_/n3 ), .a(\net237[10] ) );
    inv_1 \U14_5_/U4  ( .x(\U14_5_/n4 ), .a(\net246[10] ) );
    inv_1 \U14_5_/U5  ( .x(\net212[10] ), .a(\U14_5_/n5 ) );
    and4_1 \U14_6_/U16  ( .x(\U14_6_/n5 ), .a(\U14_6_/n1 ), .b(\U14_6_/n2 ), 
        .c(\U14_6_/n3 ), .d(\U14_6_/n4 ) );
    inv_1 \U14_6_/U1  ( .x(\U14_6_/n1 ), .a(\net231[9] ) );
    inv_1 \U14_6_/U2  ( .x(\U14_6_/n2 ), .a(\net222[9] ) );
    inv_1 \U14_6_/U3  ( .x(\U14_6_/n3 ), .a(\net237[9] ) );
    inv_1 \U14_6_/U4  ( .x(\U14_6_/n4 ), .a(\net246[9] ) );
    inv_1 \U14_6_/U5  ( .x(\net212[9] ), .a(\U14_6_/n5 ) );
    and4_1 \U14_7_/U16  ( .x(\U14_7_/n5 ), .a(\U14_7_/n1 ), .b(\U14_7_/n2 ), 
        .c(\U14_7_/n3 ), .d(\U14_7_/n4 ) );
    inv_1 \U14_7_/U1  ( .x(\U14_7_/n1 ), .a(\net231[8] ) );
    inv_1 \U14_7_/U2  ( .x(\U14_7_/n2 ), .a(\net222[8] ) );
    inv_1 \U14_7_/U3  ( .x(\U14_7_/n3 ), .a(\net237[8] ) );
    inv_1 \U14_7_/U4  ( .x(\U14_7_/n4 ), .a(\net246[8] ) );
    inv_1 \U14_7_/U5  ( .x(\net212[8] ), .a(\U14_7_/n5 ) );
    and4_1 \U14_8_/U16  ( .x(\U14_8_/n5 ), .a(\U14_8_/n1 ), .b(\U14_8_/n2 ), 
        .c(\U14_8_/n3 ), .d(\U14_8_/n4 ) );
    inv_1 \U14_8_/U1  ( .x(\U14_8_/n1 ), .a(\net231[7] ) );
    inv_1 \U14_8_/U2  ( .x(\U14_8_/n2 ), .a(\net222[7] ) );
    inv_1 \U14_8_/U3  ( .x(\U14_8_/n3 ), .a(\net237[7] ) );
    inv_1 \U14_8_/U4  ( .x(\U14_8_/n4 ), .a(\net246[7] ) );
    inv_1 \U14_8_/U5  ( .x(\net212[7] ), .a(\U14_8_/n5 ) );
    and4_1 \U14_9_/U16  ( .x(\U14_9_/n5 ), .a(\U14_9_/n1 ), .b(\U14_9_/n2 ), 
        .c(\U14_9_/n3 ), .d(\U14_9_/n4 ) );
    inv_1 \U14_9_/U1  ( .x(\U14_9_/n1 ), .a(\net231[6] ) );
    inv_1 \U14_9_/U2  ( .x(\U14_9_/n2 ), .a(\net222[6] ) );
    inv_1 \U14_9_/U3  ( .x(\U14_9_/n3 ), .a(\net237[6] ) );
    inv_1 \U14_9_/U4  ( .x(\U14_9_/n4 ), .a(\net246[6] ) );
    inv_1 \U14_9_/U5  ( .x(\net212[6] ), .a(\U14_9_/n5 ) );
    and4_1 \U14_10_/U16  ( .x(\U14_10_/n5 ), .a(\U14_10_/n1 ), .b(\U14_10_/n2 
        ), .c(\U14_10_/n3 ), .d(\U14_10_/n4 ) );
    inv_1 \U14_10_/U1  ( .x(\U14_10_/n1 ), .a(\net231[5] ) );
    inv_1 \U14_10_/U2  ( .x(\U14_10_/n2 ), .a(\net222[5] ) );
    inv_1 \U14_10_/U3  ( .x(\U14_10_/n3 ), .a(\net237[5] ) );
    inv_1 \U14_10_/U4  ( .x(\U14_10_/n4 ), .a(\net246[5] ) );
    inv_1 \U14_10_/U5  ( .x(\net212[5] ), .a(\U14_10_/n5 ) );
    inv_1 \U14_11_/U1  ( .x(\U14_11_/n1 ), .a(\net231[4] ) );
    inv_1 \U14_11_/U2  ( .x(\U14_11_/n2 ), .a(\net222[4] ) );
    inv_1 \U14_11_/U4  ( .x(\U14_11_/n4 ), .a(\net246[4] ) );
    inv_1 \U14_11_/U5  ( .x(\net212[4] ), .a(\U14_11_/n5 ) );
    inv_1 \U14_12_/U1  ( .x(\U14_12_/n1 ), .a(\net231[3] ) );
    inv_1 \U14_12_/U2  ( .x(\U14_12_/n2 ), .a(\net222[3] ) );
    inv_1 \U14_12_/U4  ( .x(\U14_12_/n4 ), .a(\net246[3] ) );
    inv_1 \U14_12_/U5  ( .x(\net212[3] ), .a(\U14_12_/n5 ) );
    and4_1 \U14_13_/U16  ( .x(\U14_13_/n5 ), .a(\U14_13_/n1 ), .b(\U14_13_/n2 
        ), .c(\U14_13_/n3 ), .d(\U14_13_/n4 ) );
    inv_1 \U14_13_/U1  ( .x(\U14_13_/n1 ), .a(\net231[2] ) );
    inv_1 \U14_13_/U2  ( .x(\U14_13_/n2 ), .a(\net222[2] ) );
    inv_1 \U14_13_/U3  ( .x(\U14_13_/n3 ), .a(\net237[2] ) );
    inv_1 \U14_13_/U4  ( .x(\U14_13_/n4 ), .a(\net246[2] ) );
    inv_1 \U14_13_/U5  ( .x(\net212[2] ), .a(\U14_13_/n5 ) );
    and4_1 \U14_14_/U16  ( .x(\U14_14_/n5 ), .a(\U14_14_/n1 ), .b(\U14_14_/n2 
        ), .c(\U14_14_/n3 ), .d(\U14_14_/n4 ) );
    inv_1 \U14_14_/U1  ( .x(\U14_14_/n1 ), .a(\net231[1] ) );
    inv_1 \U14_14_/U2  ( .x(\U14_14_/n2 ), .a(\net222[1] ) );
    inv_1 \U14_14_/U3  ( .x(\U14_14_/n3 ), .a(\net237[1] ) );
    inv_1 \U14_14_/U4  ( .x(\U14_14_/n4 ), .a(\net246[1] ) );
    inv_1 \U14_14_/U5  ( .x(\net212[1] ), .a(\U14_14_/n5 ) );
    and4_1 \U14_15_/U16  ( .x(\U14_15_/n5 ), .a(\U14_15_/n1 ), .b(\U14_15_/n2 
        ), .c(\U14_15_/n3 ), .d(\U14_15_/n4 ) );
    inv_1 \U14_15_/U1  ( .x(\U14_15_/n1 ), .a(\net231[0] ) );
    inv_1 \U14_15_/U2  ( .x(\U14_15_/n2 ), .a(\net222[0] ) );
    inv_1 \U14_15_/U3  ( .x(\U14_15_/n3 ), .a(\net237[0] ) );
    inv_1 \U14_15_/U4  ( .x(\U14_15_/n4 ), .a(\net246[0] ) );
    inv_1 \U14_15_/U5  ( .x(\net212[0] ), .a(\U14_15_/n5 ) );
    and4_1 \U91_0_/U16  ( .x(\U91_0_/n5 ), .a(\U91_0_/n1 ), .b(\U91_0_/n2 ), 
        .c(\U91_0_/n3 ), .d(\U91_0_/n4 ) );
    inv_1 \U91_0_/U1  ( .x(\U91_0_/n1 ), .a(\net219[15] ) );
    inv_1 \U91_0_/U2  ( .x(\U91_0_/n2 ), .a(\net243[15] ) );
    inv_1 \U91_0_/U3  ( .x(\U91_0_/n3 ), .a(\net240[15] ) );
    inv_1 \U91_0_/U4  ( .x(\U91_0_/n4 ), .a(\net228[15] ) );
    inv_1 \U91_0_/U5  ( .x(\net207[15] ), .a(\U91_0_/n5 ) );
    and4_1 \U91_1_/U16  ( .x(\U91_1_/n5 ), .a(\U91_1_/n1 ), .b(\U91_1_/n2 ), 
        .c(\U91_1_/n3 ), .d(\U91_1_/n4 ) );
    inv_1 \U91_1_/U1  ( .x(\U91_1_/n1 ), .a(\net219[14] ) );
    inv_1 \U91_1_/U2  ( .x(\U91_1_/n2 ), .a(\net243[14] ) );
    inv_1 \U91_1_/U3  ( .x(\U91_1_/n3 ), .a(\net240[14] ) );
    inv_1 \U91_1_/U4  ( .x(\U91_1_/n4 ), .a(\net228[14] ) );
    inv_1 \U91_1_/U5  ( .x(\net207[14] ), .a(\U91_1_/n5 ) );
    and4_1 \U91_2_/U16  ( .x(\U91_2_/n5 ), .a(\U91_2_/n1 ), .b(\U91_2_/n2 ), 
        .c(\U91_2_/n3 ), .d(\U91_2_/n4 ) );
    inv_1 \U91_2_/U1  ( .x(\U91_2_/n1 ), .a(\net219[13] ) );
    inv_1 \U91_2_/U2  ( .x(\U91_2_/n2 ), .a(\net243[13] ) );
    inv_1 \U91_2_/U3  ( .x(\U91_2_/n3 ), .a(\net240[13] ) );
    inv_1 \U91_2_/U4  ( .x(\U91_2_/n4 ), .a(\net228[13] ) );
    inv_1 \U91_2_/U5  ( .x(\net207[13] ), .a(\U91_2_/n5 ) );
    and4_1 \U91_3_/U16  ( .x(\U91_3_/n5 ), .a(\U91_3_/n1 ), .b(\U91_3_/n2 ), 
        .c(\U91_3_/n3 ), .d(\U91_3_/n4 ) );
    inv_1 \U91_3_/U1  ( .x(\U91_3_/n1 ), .a(\net219[12] ) );
    inv_1 \U91_3_/U2  ( .x(\U91_3_/n2 ), .a(\net243[12] ) );
    inv_1 \U91_3_/U3  ( .x(\U91_3_/n3 ), .a(\net240[12] ) );
    inv_1 \U91_3_/U4  ( .x(\U91_3_/n4 ), .a(\net228[12] ) );
    inv_1 \U91_3_/U5  ( .x(\net207[12] ), .a(\U91_3_/n5 ) );
    and4_1 \U91_4_/U16  ( .x(\U91_4_/n5 ), .a(\U91_4_/n1 ), .b(\U91_4_/n2 ), 
        .c(\U91_4_/n3 ), .d(\U91_4_/n4 ) );
    inv_1 \U91_4_/U1  ( .x(\U91_4_/n1 ), .a(\net219[11] ) );
    inv_1 \U91_4_/U2  ( .x(\U91_4_/n2 ), .a(\net243[11] ) );
    inv_1 \U91_4_/U3  ( .x(\U91_4_/n3 ), .a(\net240[11] ) );
    inv_1 \U91_4_/U4  ( .x(\U91_4_/n4 ), .a(\net228[11] ) );
    inv_1 \U91_4_/U5  ( .x(\net207[11] ), .a(\U91_4_/n5 ) );
    and4_1 \U91_5_/U16  ( .x(\U91_5_/n5 ), .a(\U91_5_/n1 ), .b(\U91_5_/n2 ), 
        .c(\U91_5_/n3 ), .d(\U91_5_/n4 ) );
    inv_1 \U91_5_/U1  ( .x(\U91_5_/n1 ), .a(\net219[10] ) );
    inv_1 \U91_5_/U2  ( .x(\U91_5_/n2 ), .a(\net243[10] ) );
    inv_1 \U91_5_/U3  ( .x(\U91_5_/n3 ), .a(\net240[10] ) );
    inv_1 \U91_5_/U4  ( .x(\U91_5_/n4 ), .a(\net228[10] ) );
    inv_1 \U91_5_/U5  ( .x(\net207[10] ), .a(\U91_5_/n5 ) );
    and4_1 \U91_6_/U16  ( .x(\U91_6_/n5 ), .a(\U91_6_/n1 ), .b(\U91_6_/n2 ), 
        .c(\U91_6_/n3 ), .d(\U91_6_/n4 ) );
    inv_1 \U91_6_/U1  ( .x(\U91_6_/n1 ), .a(\net219[9] ) );
    inv_1 \U91_6_/U2  ( .x(\U91_6_/n2 ), .a(\net243[9] ) );
    inv_1 \U91_6_/U3  ( .x(\U91_6_/n3 ), .a(\net240[9] ) );
    inv_1 \U91_6_/U4  ( .x(\U91_6_/n4 ), .a(\net228[9] ) );
    inv_1 \U91_6_/U5  ( .x(\net207[9] ), .a(\U91_6_/n5 ) );
    and4_1 \U91_7_/U16  ( .x(\U91_7_/n5 ), .a(\U91_7_/n1 ), .b(\U91_7_/n2 ), 
        .c(\U91_7_/n3 ), .d(\U91_7_/n4 ) );
    inv_1 \U91_7_/U1  ( .x(\U91_7_/n1 ), .a(\net219[8] ) );
    inv_1 \U91_7_/U2  ( .x(\U91_7_/n2 ), .a(\net243[8] ) );
    inv_1 \U91_7_/U3  ( .x(\U91_7_/n3 ), .a(\net240[8] ) );
    inv_1 \U91_7_/U4  ( .x(\U91_7_/n4 ), .a(\net228[8] ) );
    inv_1 \U91_7_/U5  ( .x(\net207[8] ), .a(\U91_7_/n5 ) );
    and4_1 \U91_8_/U16  ( .x(\U91_8_/n5 ), .a(\U91_8_/n1 ), .b(\U91_8_/n2 ), 
        .c(\U91_8_/n3 ), .d(\U91_8_/n4 ) );
    inv_1 \U91_8_/U1  ( .x(\U91_8_/n1 ), .a(\net219[7] ) );
    inv_1 \U91_8_/U2  ( .x(\U91_8_/n2 ), .a(\net243[7] ) );
    inv_1 \U91_8_/U3  ( .x(\U91_8_/n3 ), .a(\net240[7] ) );
    inv_1 \U91_8_/U4  ( .x(\U91_8_/n4 ), .a(\net228[7] ) );
    inv_1 \U91_8_/U5  ( .x(\net207[7] ), .a(\U91_8_/n5 ) );
    and4_1 \U91_9_/U16  ( .x(\U91_9_/n5 ), .a(\U91_9_/n1 ), .b(\U91_9_/n2 ), 
        .c(\U91_9_/n3 ), .d(\U91_9_/n4 ) );
    inv_1 \U91_9_/U1  ( .x(\U91_9_/n1 ), .a(\net219[6] ) );
    inv_1 \U91_9_/U2  ( .x(\U91_9_/n2 ), .a(\net243[6] ) );
    inv_1 \U91_9_/U3  ( .x(\U91_9_/n3 ), .a(\net240[6] ) );
    inv_1 \U91_9_/U4  ( .x(\U91_9_/n4 ), .a(\net228[6] ) );
    inv_1 \U91_9_/U5  ( .x(\net207[6] ), .a(\U91_9_/n5 ) );
    and4_1 \U91_10_/U16  ( .x(\U91_10_/n5 ), .a(\U91_10_/n1 ), .b(\U91_10_/n2 
        ), .c(\U91_10_/n3 ), .d(\U91_10_/n4 ) );
    inv_1 \U91_10_/U1  ( .x(\U91_10_/n1 ), .a(\net219[5] ) );
    inv_1 \U91_10_/U2  ( .x(\U91_10_/n2 ), .a(\net243[5] ) );
    inv_1 \U91_10_/U3  ( .x(\U91_10_/n3 ), .a(\net240[5] ) );
    inv_1 \U91_10_/U4  ( .x(\U91_10_/n4 ), .a(\net228[5] ) );
    inv_1 \U91_10_/U5  ( .x(\net207[5] ), .a(\U91_10_/n5 ) );
    and4_1 \U91_11_/U16  ( .x(\U91_11_/n5 ), .a(\U91_11_/n1 ), .b(\U91_11_/n2 
        ), .c(\U91_11_/n3 ), .d(\U91_11_/n4 ) );
    inv_1 \U91_11_/U1  ( .x(\U91_11_/n1 ), .a(\net219[4] ) );
    inv_1 \U91_11_/U2  ( .x(\U91_11_/n2 ), .a(\net243[4] ) );
    inv_1 \U91_11_/U3  ( .x(\U91_11_/n3 ), .a(\net240[4] ) );
    inv_1 \U91_11_/U4  ( .x(\U91_11_/n4 ), .a(\net228[4] ) );
    inv_1 \U91_11_/U5  ( .x(\net207[4] ), .a(\U91_11_/n5 ) );
    and4_1 \U91_12_/U16  ( .x(\U91_12_/n5 ), .a(\U91_12_/n1 ), .b(\U91_12_/n2 
        ), .c(\U91_12_/n3 ), .d(\U91_12_/n4 ) );
    inv_1 \U91_12_/U1  ( .x(\U91_12_/n1 ), .a(\net219[3] ) );
    inv_1 \U91_12_/U2  ( .x(\U91_12_/n2 ), .a(\net243[3] ) );
    inv_1 \U91_12_/U3  ( .x(\U91_12_/n3 ), .a(\net240[3] ) );
    inv_1 \U91_12_/U4  ( .x(\U91_12_/n4 ), .a(\net228[3] ) );
    inv_1 \U91_12_/U5  ( .x(\net207[3] ), .a(\U91_12_/n5 ) );
    and4_1 \U91_13_/U16  ( .x(\U91_13_/n5 ), .a(\U91_13_/n1 ), .b(\U91_13_/n2 
        ), .c(\U91_13_/n3 ), .d(\U91_13_/n4 ) );
    inv_1 \U91_13_/U1  ( .x(\U91_13_/n1 ), .a(\net219[2] ) );
    inv_1 \U91_13_/U2  ( .x(\U91_13_/n2 ), .a(\net243[2] ) );
    inv_1 \U91_13_/U3  ( .x(\U91_13_/n3 ), .a(\net240[2] ) );
    inv_1 \U91_13_/U4  ( .x(\U91_13_/n4 ), .a(\net228[2] ) );
    inv_1 \U91_13_/U5  ( .x(\net207[2] ), .a(\U91_13_/n5 ) );
    and4_1 \U91_14_/U16  ( .x(\U91_14_/n5 ), .a(\U91_14_/n1 ), .b(\U91_14_/n2 
        ), .c(\U91_14_/n3 ), .d(\U91_14_/n4 ) );
    inv_1 \U91_14_/U1  ( .x(\U91_14_/n1 ), .a(\net219[1] ) );
    inv_1 \U91_14_/U2  ( .x(\U91_14_/n2 ), .a(\net243[1] ) );
    inv_1 \U91_14_/U3  ( .x(\U91_14_/n3 ), .a(\net240[1] ) );
    inv_1 \U91_14_/U4  ( .x(\U91_14_/n4 ), .a(\net228[1] ) );
    inv_1 \U91_14_/U5  ( .x(\net207[1] ), .a(\U91_14_/n5 ) );
    and4_1 \U91_15_/U16  ( .x(\U91_15_/n5 ), .a(\U91_15_/n1 ), .b(\U91_15_/n2 
        ), .c(\U91_15_/n3 ), .d(\U91_15_/n4 ) );
    inv_1 \U91_15_/U1  ( .x(\U91_15_/n1 ), .a(\net219[0] ) );
    inv_1 \U91_15_/U2  ( .x(\U91_15_/n2 ), .a(\net243[0] ) );
    inv_1 \U91_15_/U3  ( .x(\U91_15_/n3 ), .a(\net240[0] ) );
    inv_1 \U91_15_/U4  ( .x(\U91_15_/n4 ), .a(\net228[0] ) );
    inv_1 \U91_15_/U5  ( .x(\net207[0] ), .a(\U91_15_/n5 ) );
    or3_2 \U93_0_/U12  ( .x(chainl[0]), .a(\net207[15] ), .b(\net217[15] ), 
        .c(\net212[15] ) );
    or3_2 \U93_1_/U12  ( .x(chainl[1]), .a(\net207[14] ), .b(\net217[14] ), 
        .c(\net212[14] ) );
    or3_2 \U93_2_/U12  ( .x(chainl[2]), .a(\net207[13] ), .b(\net217[13] ), 
        .c(\net212[13] ) );
    or3_2 \U93_3_/U12  ( .x(chainl[3]), .a(\net207[12] ), .b(\net217[12] ), 
        .c(\net212[12] ) );
    or3_2 \U93_4_/U12  ( .x(chainl[4]), .a(\net207[11] ), .b(\net217[11] ), 
        .c(\net212[11] ) );
    or3_2 \U93_5_/U12  ( .x(chainl[5]), .a(\net207[10] ), .b(\net217[10] ), 
        .c(\net212[10] ) );
    or3_2 \U93_6_/U12  ( .x(chainl[6]), .a(\net207[9] ), .b(\net217[9] ), .c(
        \net212[9] ) );
    or3_2 \U93_7_/U12  ( .x(chainl[7]), .a(\net207[8] ), .b(\net217[8] ), .c(
        \net212[8] ) );
    or3_2 \U93_8_/U12  ( .x(chainh[0]), .a(\net207[7] ), .b(\net217[7] ), .c(
        \net212[7] ) );
    or3_2 \U93_9_/U12  ( .x(chainh[1]), .a(\net207[6] ), .b(\net217[6] ), .c(
        \net212[6] ) );
    or3_2 \U93_10_/U12  ( .x(chainh[2]), .a(\net207[5] ), .b(\net217[5] ), .c(
        \net212[5] ) );
    or3_2 \U93_11_/U12  ( .x(chainh[3]), .a(\net207[4] ), .b(\net217[4] ), .c(
        \net212[4] ) );
    or3_2 \U93_12_/U12  ( .x(chainh[4]), .a(\net207[3] ), .b(\net217[3] ), .c(
        \net212[3] ) );
    or3_2 \U93_13_/U12  ( .x(chainh[5]), .a(\net207[2] ), .b(\net217[2] ), .c(
        \net212[2] ) );
    or3_2 \U93_14_/U12  ( .x(chainh[6]), .a(\net207[1] ), .b(\net217[1] ), .c(
        \net212[1] ) );
    or3_2 \U93_15_/U12  ( .x(chainh[7]), .a(\net207[0] ), .b(\net217[0] ), .c(
        \net212[0] ) );
    inv_1 \U152/U3  ( .x(net198), .a(sendreq) );
    ao23_1 \U158/U19/U21/U1/U1  ( .x(net131), .a(net132), .b(net131), .c(
        net132), .d(rnw[1]), .e(rnw[1]) );
    ao23_1 \U157/U19/U21/U1/U1  ( .x(net176), .a(net132), .b(net176), .c(
        net132), .d(rnw[0]), .e(rnw[0]) );
    ao222_1 \U123/U18/U1/U1  ( .x(net136), .a(net185), .b(net187), .c(net185), 
        .d(net136), .e(net187), .f(net136) );
    aoi21_1 \U151/U30/U1/U1  ( .x(\hdr[4] ), .a(\U151/Z ), .b(net138), .c(
        net198) );
    inv_1 \U151/U30/U1/U2  ( .x(\U151/Z ), .a(\hdr[4] ) );
    nor3_1 \U148/U21/Unr  ( .x(\U148/U21/nr ), .a(net191), .b(net136), .c(
        net293) );
    nand3_1 \U148/U21/Und  ( .x(\U148/U21/nd ), .a(net191), .b(net136), .c(
        net293) );
    oa21_1 \U148/U21/U1  ( .x(\U148/U21/n2 ), .a(\U148/U21/n2 ), .b(
        \U148/U21/nr ), .c(\U148/U21/nd ) );
    inv_1 \U148/U21/U3  ( .x(ack), .a(\U148/U21/n2 ) );
    buf_3 U1 ( .x(n1), .a(net138) );
    buf_3 U2 ( .x(net138), .a(nia) );
    buf_3 U3 ( .x(net269), .a(net146) );
    buf_3 U4 ( .x(net255), .a(\bs[5] ) );
    buf_3 U5 ( .x(net267), .a(\bs[6] ) );
    buf_3 U6 ( .x(net253), .a(\bs[2] ) );
    buf_3 U7 ( .x(net249), .a(\bs[8] ) );
    buf_3 U8 ( .x(net263), .a(\bs[7] ) );
    buf_3 U9 ( .x(net259), .a(\bs[3] ) );
    buf_3 U10 ( .x(net251), .a(\bs[4] ) );
    buf_3 U11 ( .x(net261), .a(\bs[1] ) );
    buf_3 U12 ( .x(net265), .a(\bs[0] ) );
    and2_1 U13 ( .x(\U40_2_/n5 ), .a(\U40_2_/n3 ), .b(\U40_2_/n4 ) );
    and2_1 U14 ( .x(\U40_1_/n5 ), .a(\U40_1_/n3 ), .b(\U40_1_/n4 ) );
    and2_1 U15 ( .x(\U40_9_/n5 ), .a(\U40_9_/n3 ), .b(\U40_9_/n4 ) );
    and2_1 U16 ( .x(\U40_8_/n5 ), .a(\U40_8_/n3 ), .b(\U40_8_/n4 ) );
    and2_1 U17 ( .x(\U40_13_/n5 ), .a(\U40_13_/n3 ), .b(\U40_13_/n4 ) );
    and2_1 U18 ( .x(\U40_0_/n5 ), .a(\U40_0_/n3 ), .b(\U40_0_/n4 ) );
    and2_1 U19 ( .x(\U40_5_/n5 ), .a(\U40_5_/n3 ), .b(\U40_5_/n4 ) );
    and2_1 U20 ( .x(\U40_4_/n5 ), .a(\U40_4_/n3 ), .b(\U40_4_/n4 ) );
    and3_1 U21 ( .x(\U14_12_/n5 ), .a(\U14_12_/n2 ), .b(\U14_12_/n4 ), .c(
        \U14_12_/n1 ) );
    and2_1 U22 ( .x(\U40_12_/n5 ), .a(\U40_12_/n3 ), .b(\U40_12_/n4 ) );
    and2_1 U23 ( .x(\U40_3_/n5 ), .a(\U40_3_/n3 ), .b(\U40_3_/n4 ) );
    and3_1 U24 ( .x(\U14_11_/n5 ), .a(\U14_11_/n2 ), .b(\U14_11_/n4 ), .c(
        \U14_11_/n1 ) );
    and2_1 U25 ( .x(\U40_11_/n5 ), .a(\U40_11_/n3 ), .b(\U40_11_/n4 ) );
    and2_1 U26 ( .x(\U40_10_/n5 ), .a(\U40_10_/n3 ), .b(\U40_10_/n4 ) );
    and2_1 U27 ( .x(\U40_15_/n5 ), .a(\U40_15_/n3 ), .b(\U40_15_/n4 ) );
    and2_1 U28 ( .x(\U40_7_/n5 ), .a(\U40_7_/n3 ), .b(\U40_7_/n4 ) );
    and2_1 U29 ( .x(\U40_6_/n5 ), .a(\U40_6_/n3 ), .b(\U40_6_/n4 ) );
    and2_1 U30 ( .x(\U40_14_/n5 ), .a(\U40_14_/n3 ), .b(\U40_14_/n4 ) );
endmodule


module chain_ic_ctrl_2 ( ack, candefer, eop, nstatack, pltxreq, routetxreq, 
    tok_ack, accept, candefer_ack, defer, eopack, lock, nReset, pltxack, 
    routetxack, tok_err, tok_ok );
input  [1:0] candefer_ack;
input  [1:0] lock;
input  accept, defer, eopack, nReset, pltxack, routetxack, tok_err, tok_ok;
output ack, candefer, eop, nstatack, pltxreq, routetxreq, tok_ack;
    wire \locked[1] , \locked[0] , net21, net12, net20, net16, net10, net7, 
        net6, retry, net27, txnodefer, net13, txunlocked, net5, txmaydefer, 
        txdone, net8, txlocked, net29, net2, net4, lockcleared, net28, net18, 
        net22, net14, net9, net24, net19, net31, net11, net30, net17, net3, 
        reset, net26, nlclear, lwrite, net15, net23, net25, \U249/n5 , 
        \U249/n1 , \U249/n2 , \U249/n3 , \U249/n4 , \U286/U28/U1/clr , 
        \U286/U28/U1/set , \U285/U28/U1/clr , \U285/U28/U1/set , 
        \U262/U25/U1/clr , \U262/U25/U1/ob , \U284/U25/U1/clr , 
        \U284/U25/U1/ob , \U283/U25/U1/clr , \U283/U25/U1/ob , \U288/Z , 
        \U289/Z , \U287/Z , \U149/nr , \U149/nd , \U149/n2 , \U160/acb , 
        \U160/U1/Z , \U136/nlsense , \U136/nulsense , \U136/nwh , \U136/nwl , 
        \U136/nclear_latch , n1, n2;
    nand2_1 \U146/U5  ( .x(candefer), .a(net23), .b(net25) );
    or2_1 \U277/U12  ( .x(net6), .a(net19), .b(net9) );
    or2_1 \U264/U12  ( .x(retry), .a(net31), .b(net24) );
    or2_1 \U259/U12  ( .x(net28), .a(net27), .b(net7) );
    or2_1 \U140/U12  ( .x(net18), .a(net13), .b(net8) );
    or2_1 \U148/U12  ( .x(net11), .a(net15), .b(routetxack) );
    and4_1 \U249/U16  ( .x(\U249/n5 ), .a(\U249/n1 ), .b(\U249/n2 ), .c(
        \U249/n3 ), .d(\U249/n4 ) );
    inv_1 \U249/U1  ( .x(\U249/n1 ), .a(txnodefer) );
    inv_1 \U249/U2  ( .x(\U249/n2 ), .a(net16) );
    inv_1 \U249/U3  ( .x(\U249/n3 ), .a(net9) );
    inv_1 \U249/U4  ( .x(\U249/n4 ), .a(net19) );
    inv_1 \U249/U5  ( .x(ack), .a(\U249/n5 ) );
    nor3_2 \U40/U16  ( .x(nstatack), .a(net16), .b(reset), .c(retry) );
    nor3_2 \U275/U16  ( .x(net17), .a(net29), .b(reset), .c(tok_ack) );
    buf_3 \U290/U8  ( .x(net12), .a(txmaydefer) );
    nor2_1 \U154/U5  ( .x(nlclear), .a(net4), .b(net31) );
    or2_2 \U274/U12  ( .x(pltxreq), .a(net22), .b(net14) );
    or3_1 \U260/U12  ( .x(eop), .a(net31), .b(txlocked), .c(net4) );
    inv_1 \U147/U3  ( .x(net3), .a(net29) );
    inv_1 \U174/U3  ( .x(reset), .a(nReset) );
    aoai211_1 \U286/U28/U1/U1  ( .x(\U286/U28/U1/clr ), .a(net3), .b(n1), .c(
        net17), .d(net22) );
    nand3_1 \U286/U28/U1/U2  ( .x(\U286/U28/U1/set ), .a(net17), .b(net3), .c(
        n1) );
    nand2_2 \U286/U28/U1/U3  ( .x(net22), .a(\U286/U28/U1/clr ), .b(
        \U286/U28/U1/set ) );
    aoai211_1 \U285/U28/U1/U1  ( .x(\U285/U28/U1/clr ), .a(net3), .b(n2), .c(
        net17), .d(net14) );
    nand3_1 \U285/U28/U1/U2  ( .x(\U285/U28/U1/set ), .a(net17), .b(net3), .c(
        n2) );
    nand2_2 \U285/U28/U1/U3  ( .x(net14), .a(\U285/U28/U1/clr ), .b(
        \U285/U28/U1/set ) );
    ao222_1 \U254/U18/U1/U1  ( .x(net31), .a(defer), .b(txunlocked), .c(defer), 
        .d(net31), .e(txunlocked), .f(net31) );
    ao222_1 \U252/U18/U1/U1  ( .x(net19), .a(tok_err), .b(net12), .c(tok_err), 
        .d(net19), .e(net12), .f(net19) );
    ao222_1 \U276/U18/U1/U1  ( .x(net24), .a(txlocked), .b(defer), .c(txlocked
        ), .d(net24), .e(defer), .f(net24) );
    ao222_1 \U251/U18/U1/U1  ( .x(net9), .a(tok_ok), .b(net12), .c(tok_ok), 
        .d(net9), .e(net12), .f(net9) );
    ao222_1 \U235/U18/U1/U1  ( .x(tok_ack), .a(ack), .b(net2), .c(ack), .d(
        tok_ack), .e(net2), .f(tok_ack) );
    ao222_1 \U247/U18/U1/U1  ( .x(txnodefer), .a(txdone), .b(candefer_ack[0]), 
        .c(txdone), .d(txnodefer), .e(candefer_ack[0]), .f(txnodefer) );
    ao222_2 \U246/U19/U1/U1  ( .x(txlocked), .a(net14), .b(txdone), .c(net14), 
        .d(txlocked), .e(txdone), .f(txlocked) );
    ao222_2 \U245/U19/U1/U1  ( .x(txunlocked), .a(txdone), .b(net22), .c(
        txdone), .d(txunlocked), .e(net22), .f(txunlocked) );
    ao222_1 \U269/U18/U1/U1  ( .x(net2), .a(net28), .b(net18), .c(net28), .d(
        net2), .e(net18), .f(net2) );
    ao222_1 \U268/U18/U1/U1  ( .x(net5), .a(eopack), .b(lockcleared), .c(
        eopack), .d(net5), .e(lockcleared), .f(net5) );
    ao222_1 \U256/U18/U1/U1  ( .x(net4), .a(tok_err), .b(txunlocked), .c(
        tok_err), .d(net4), .e(txunlocked), .f(net4) );
    ao222_1 \U175/U18/U1/U1  ( .x(net29), .a(net2), .b(retry), .c(net2), .d(
        net29), .e(retry), .f(net29) );
    ao222_1 \U255/U18/U1/U1  ( .x(net8), .a(txlocked), .b(eopack), .c(txlocked
        ), .d(net8), .e(eopack), .f(net8) );
    ao222_2 \U248/U19/U1/U1  ( .x(txmaydefer), .a(candefer_ack[1]), .b(txdone), 
        .c(candefer_ack[1]), .d(txmaydefer), .e(txdone), .f(txmaydefer) );
    ao222_2 \U250/U19/U1/U1  ( .x(net16), .a(accept), .b(net12), .c(accept), 
        .d(net16), .e(net12), .f(net16) );
    oa31_1 \U262/U25/U1/Uclr  ( .x(\U262/U25/U1/clr ), .a(txunlocked), .b(net5
        ), .c(tok_ok), .d(net13) );
    oaoi211_1 \U262/U25/U1/Uaoi  ( .x(\U262/U25/U1/ob ), .a(net5), .b(tok_ok), 
        .c(txunlocked), .d(\U262/U25/U1/clr ) );
    inv_2 \U262/U25/U1/Ui  ( .x(net13), .a(\U262/U25/U1/ob ) );
    oa31_1 \U284/U25/U1/Uclr  ( .x(\U284/U25/U1/clr ), .a(txnodefer), .b(
        tok_ok), .c(tok_err), .d(net27) );
    oaoi211_1 \U284/U25/U1/Uaoi  ( .x(\U284/U25/U1/ob ), .a(tok_ok), .b(
        tok_err), .c(txnodefer), .d(\U284/U25/U1/clr ) );
    inv_2 \U284/U25/U1/Ui  ( .x(net27), .a(\U284/U25/U1/ob ) );
    oa31_1 \U283/U25/U1/Uclr  ( .x(\U283/U25/U1/clr ), .a(net10), .b(net6), 
        .c(retry), .d(net7) );
    oaoi211_1 \U283/U25/U1/Uaoi  ( .x(\U283/U25/U1/ob ), .a(net6), .b(retry), 
        .c(net10), .d(\U283/U25/U1/clr ) );
    inv_2 \U283/U25/U1/Ui  ( .x(net7), .a(\U283/U25/U1/ob ) );
    aoi21_1 \U289/U30/U1/U1  ( .x(net20), .a(\U289/Z ), .b(net16), .c(net12)
         );
    inv_1 \U289/U30/U1/U2  ( .x(\U289/Z ), .a(net20) );
    aoi21_1 \U287/U30/U1/U1  ( .x(net21), .a(\U287/Z ), .b(accept), .c(net12)
         );
    inv_1 \U287/U30/U1/U2  ( .x(\U287/Z ), .a(net21) );
    aoi222_1 \U288/U30/U1  ( .x(net10), .a(net20), .b(net21), .c(net20), .d(
        \U288/Z ), .e(net21), .f(\U288/Z ) );
    inv_1 \U288/U30/Uinv  ( .x(\U288/Z ), .a(net10) );
    nor3_1 \U149/Unr  ( .x(\U149/nr ), .a(pltxack), .b(net11), .c(net30) );
    nand3_1 \U149/Und  ( .x(\U149/nd ), .a(pltxack), .b(net11), .c(net30) );
    oa21_1 \U149/U1  ( .x(\U149/n2 ), .a(\U149/n2 ), .b(\U149/nr ), .c(
        \U149/nd ) );
    inv_2 \U149/U3  ( .x(txdone), .a(\U149/n2 ) );
    inv_1 \U133/U618/U3  ( .x(net23), .a(net15) );
    inv_1 \U133/U617/U3  ( .x(net25), .a(routetxreq) );
    ao23_1 \U133/U616/U21/U1/U1  ( .x(routetxreq), .a(pltxreq), .b(routetxreq), 
        .c(pltxreq), .d(\locked[0] ), .e(net23) );
    ao23_1 \U133/U615/U21/U1/U1  ( .x(net15), .a(pltxreq), .b(net15), .c(
        pltxreq), .d(\locked[1] ), .e(net25) );
    and2_1 \U160/U2/U8  ( .x(lwrite), .a(candefer), .b(\U160/acb ) );
    nor2_1 \U160/U3/U5  ( .x(net30), .a(\U160/acb ), .b(net26) );
    oai21_1 \U160/U1/U30/U1/U1  ( .x(\U160/acb ), .a(\U160/U1/Z ), .b(net26), 
        .c(candefer) );
    inv_1 \U160/U1/U30/U1/U2  ( .x(\U160/U1/Z ), .a(\U160/acb ) );
    nand3_2 \U136/U48/U16  ( .x(\locked[0] ), .a(\locked[1] ), .b(
        \U136/nclear_latch ), .c(\U136/nwl ) );
    nor2_0 \U136/U36/U5  ( .x(\U136/nulsense ), .a(\locked[1] ), .b(\U136/nwl 
        ) );
    nor2_0 \U136/U37/U5  ( .x(\U136/nlsense ), .a(\U136/nwh ), .b(\locked[0] )
         );
    and2_1 \U136/U76/U8  ( .x(\U136/nclear_latch ), .a(nReset), .b(nlclear) );
    nor2_1 \U136/U77/U5  ( .x(lockcleared), .a(nlclear), .b(\locked[1] ) );
    nand2_1 \U136/U14/U5  ( .x(\U136/nwl ), .a(lwrite), .b(n2) );
    nand2_1 \U136/U15/U5  ( .x(\U136/nwh ), .a(n1), .b(lwrite) );
    nand2_2 \U136/U47/U5  ( .x(\locked[1] ), .a(\U136/nwh ), .b(\locked[0] )
         );
    or2_4 \U136/U35/U12  ( .x(net26), .a(\U136/nlsense ), .b(\U136/nulsense )
         );
    buf_1 U1 ( .x(n1), .a(lock[1]) );
    buf_1 U2 ( .x(n2), .a(lock[0]) );
endmodule


module chain_irdemuxNew_2 ( err, ncback, rd, rnw, status, cbh, cbl, nReset, 
    nack, statusack );
output [1:0] err;
output [63:0] rd;
output [1:0] rnw;
output [1:0] status;
input  [7:0] cbh;
input  [7:0] cbl;
input  nReset, nack, statusack;
output ncback;
    wire n17, n18, \ncd[7] , \ncd[6] , \ncd[5] , \ncd[4] , \ncd[3] , \ncd[2] , 
        \ncd[1] , \ncd[0] , \col_h[2] , \col_h[1] , \col_h[0] , \col_l[2] , 
        \col_l[1] , \col_l[0] , \opc_l[2] , \opc_l[1] , \opc_l[0] , \opc_h[1] , 
        \opc_h[0] , pullcd, net86, net171, net168, net103, net170, bpullcd, 
        reset, net94, read_lhw, net166, net169, read, net139, net172, 
        start_receiving, net193, net167, net149, net173, pkt_normal, notify, 
        net150, write, net176, net162, pkt_done, net0187, net0208, 
        \U1697/U21/nr , \U1697/U21/nd , \U1697/U21/n2 , \U307/U21/nr , 
        \U307/U21/nd , \U307/U21/n2 , \U1664/U28/Z , \U1664/U32/Z , 
        \U1664/U29/Z , \U1664/U33/Z , \U1664/U30/Z , \U1664/U31/Z , 
        \U1664/U37/Z , \U1664/y[0] , \U1664/y[1] , \U1664/x[1] , \U1664/x[3] , 
        \U1664/x[2] , \U1664/x[0] , \U1698/nr , \U1698/nd , \U1698/n2 , 
        \I6/oh[7] , \I6/oh[6] , \I6/oh[4] , \I6/oh[3] , \I6/oh[2] , \I6/ol[7] , 
        \I6/ol[6] , \I6/ol[4] , \I6/ol[3] , \I6/drivel , \I6/driveh , 
        \I6/localcd , \I6/ncd[7] , \I6/ncd[6] , \I6/ncd[5] , \I6/ncd[4] , 
        \I6/ncd[3] , \I6/ncd[2] , \I6/ncd[1] , \I6/ncd[0] , \I6/ba , 
        \I6/latch , \I6/acb , \I6/ctrlack_internal , \I6/nlocalcd , 
        \I6/U4/U28/U1/clr , \I6/U4/U28/U1/set , \I6/U1/Z , \I6/U1664/y[0] , 
        \I6/U1664/y[1] , \I6/U1664/x[1] , \I6/U1664/x[3] , \I6/U1664/x[2] , 
        \I6/U1664/x[0] , \I6/U1664/U28/Z , \I6/U1664/U32/Z , \I6/U1664/U29/Z , 
        \I6/U1664/U33/Z , \I6/U1664/U30/Z , \I6/U1664/U31/Z , \I6/U1664/U37/Z , 
        \I6/U1669/nr , \I6/U1669/nd , \I6/U1669/n2 , \U1667/drivel , 
        \U1667/driveh , \U1667/localcd , \U1667/ncd[7] , \U1667/ncd[6] , 
        \U1667/ncd[5] , \U1667/ncd[4] , \U1667/ncd[3] , \U1667/ncd[2] , 
        \U1667/ncd[1] , \U1667/ncd[0] , \U1667/ba , \U1667/latch , \U1667/acb , 
        \U1667/ctrlack_internal , \U1667/nlocalcd , \U1667/U4/U28/U1/clr , 
        \U1667/U4/U28/U1/set , \U1667/U1/Z , \U1667/U1664/y[0] , 
        \U1667/U1664/y[1] , \U1667/U1664/x[1] , \U1667/U1664/x[3] , 
        \U1667/U1664/x[2] , \U1667/U1664/x[0] , \U1667/U1664/U28/Z , 
        \U1667/U1664/U32/Z , \U1667/U1664/U29/Z , \U1667/U1664/U33/Z , 
        \U1667/U1664/U30/Z , \U1667/U1664/U31/Z , \U1667/U1664/U37/Z , 
        \U1667/U1669/nr , \U1667/U1669/nd , \U1667/U1669/n2 , \U1650/oh[4] , 
        \U1650/oh[3] , \U1650/oh[2] , \U1650/oh[1] , \U1650/oh[0] , 
        \U1650/ol[4] , \U1650/ol[3] , \U1650/ol[2] , \U1650/ol[1] , 
        \U1650/ol[0] , \U1650/drivel , \U1650/driveh , \U1650/localcd , 
        \U1650/ncd[7] , \U1650/ncd[6] , \U1650/ncd[5] , \U1650/ncd[4] , 
        \U1650/ncd[3] , \U1650/ncd[2] , \U1650/ncd[1] , \U1650/ncd[0] , 
        \U1650/ba , \U1650/latch , \U1650/acb , \U1650/ctrlack_internal , 
        \U1650/nlocalcd , \U1650/U4/U28/U1/clr , \U1650/U4/U28/U1/set , 
        \U1650/U1/Z , \U1650/U1664/y[0] , \U1650/U1664/y[1] , 
        \U1650/U1664/x[1] , \U1650/U1664/x[3] , \U1650/U1664/x[2] , 
        \U1650/U1664/x[0] , \U1650/U1664/U28/Z , \U1650/U1664/U32/Z , 
        \U1650/U1664/U29/Z , \U1650/U1664/U33/Z , \U1650/U1664/U30/Z , 
        \U1650/U1664/U31/Z , \U1650/U1664/U37/Z , \U1650/U1669/nr , 
        \U1650/U1669/nd , \U1650/U1669/n2 , \U1666/drivel , \U1666/driveh , 
        \U1666/localcd , \U1666/ncd[7] , \U1666/ncd[6] , \U1666/ncd[5] , 
        \U1666/ncd[4] , \U1666/ncd[3] , \U1666/ncd[2] , \U1666/ncd[1] , 
        \U1666/ncd[0] , \U1666/ba , \U1666/latch , \U1666/acb , 
        \U1666/ctrlack_internal , \U1666/nlocalcd , \U1666/U4/U28/U1/clr , 
        \U1666/U4/U28/U1/set , \U1666/U1/Z , \U1666/U1664/y[0] , 
        \U1666/U1664/y[1] , \U1666/U1664/x[1] , \U1666/U1664/x[3] , 
        \U1666/U1664/x[2] , \U1666/U1664/x[0] , \U1666/U1664/U28/Z , 
        \U1666/U1664/U32/Z , \U1666/U1664/U29/Z , \U1666/U1664/U33/Z , 
        \U1666/U1664/U30/Z , \U1666/U1664/U31/Z , \U1666/U1664/U37/Z , 
        \U1666/U1669/nr , \U1666/U1669/nd , \U1666/U1669/n2 , \I1/drivel , 
        \I1/driveh , \I1/localcd , \I1/ncd[7] , \I1/ncd[6] , \I1/ncd[5] , 
        \I1/ncd[4] , \I1/ncd[3] , \I1/ncd[2] , \I1/ncd[1] , \I1/ncd[0] , 
        \I1/ba , \I1/latch , \I1/acb , \I1/ctrlack_internal , \I1/nlocalcd , 
        \I1/U4/U28/U1/clr , \I1/U4/U28/U1/set , \I1/U1/Z , \I1/U1664/y[0] , 
        \I1/U1664/y[1] , \I1/U1664/x[1] , \I1/U1664/x[3] , \I1/U1664/x[2] , 
        \I1/U1664/x[0] , \I1/U1664/U28/Z , \I1/U1664/U32/Z , \I1/U1664/U29/Z , 
        \I1/U1664/U33/Z , \I1/U1664/U30/Z , \I1/U1664/U31/Z , \I1/U1664/U37/Z , 
        \I1/U1669/nr , \I1/U1669/nd , \I1/U1669/n2 , \I2/drivel , \I2/driveh , 
        \I2/localcd , \I2/ncd[7] , \I2/ncd[6] , \I2/ncd[5] , \I2/ncd[4] , 
        \I2/ncd[3] , \I2/ncd[2] , \I2/ncd[1] , \I2/ncd[0] , \I2/ba , 
        \I2/latch , \I2/acb , \I2/ctrlack_internal , \I2/nlocalcd , 
        \I2/U4/U28/U1/clr , \I2/U4/U28/U1/set , \I2/U1/Z , \I2/U1664/y[0] , 
        \I2/U1664/y[1] , \I2/U1664/x[1] , \I2/U1664/x[3] , \I2/U1664/x[2] , 
        \I2/U1664/x[0] , \I2/U1664/U28/Z , \I2/U1664/U32/Z , \I2/U1664/U29/Z , 
        \I2/U1664/U33/Z , \I2/U1664/U30/Z , \I2/U1664/U31/Z , \I2/U1664/U37/Z , 
        \I2/U1669/nr , \I2/U1669/nd , \I2/U1669/n2 , n1, n2, n3, n4, n5, n6, 
        n7, n8, n9, n10, n11, n12, n13, n14;
    buf_1 U262 ( .x(bpullcd), .a(pullcd) );
    or2_4 \U1674/U12  ( .x(net162), .a(nack), .b(reset) );
    and2_4 \U1785/U8  ( .x(pkt_normal), .a(\opc_l[2] ), .b(\opc_l[1] ) );
    and2_4 \U1777/U8  ( .x(net150), .a(\opc_l[2] ), .b(\opc_h[1] ) );
    or3_1 \U1813/U12  ( .x(pkt_done), .a(write), .b(reset), .c(net193) );
    nor2_1 \U1651_0_/U5  ( .x(\ncd[0] ), .a(cbh[0]), .b(cbl[0]) );
    nor2_1 \U1651_1_/U5  ( .x(\ncd[1] ), .a(cbh[1]), .b(cbl[1]) );
    nor2_1 \U1651_2_/U5  ( .x(\ncd[2] ), .a(cbh[2]), .b(cbl[2]) );
    nor2_1 \U1651_3_/U5  ( .x(\ncd[3] ), .a(cbh[3]), .b(cbl[3]) );
    nor2_1 \U1651_4_/U5  ( .x(\ncd[4] ), .a(cbh[4]), .b(cbl[4]) );
    nor2_1 \U1651_5_/U5  ( .x(\ncd[5] ), .a(cbh[5]), .b(cbl[5]) );
    nor2_1 \U1651_6_/U5  ( .x(\ncd[6] ), .a(cbh[6]), .b(cbl[6]) );
    nor2_1 \U1651_7_/U5  ( .x(\ncd[7] ), .a(cbh[7]), .b(cbl[7]) );
    nor2_1 \U1812/U5  ( .x(start_receiving), .a(notify), .b(net176) );
    nor2_1 \I7/U5  ( .x(net86), .a(net172), .b(net173) );
    nor2_1 \I4/U5  ( .x(net171), .a(net169), .b(net170) );
    nor2_1 \I3/U5  ( .x(net168), .a(net166), .b(net167) );
    inv_2 \U1675/U3  ( .x(reset), .a(nReset) );
    nand3_2 \U193/U16  ( .x(ncback), .a(net86), .b(net171), .c(net168) );
    ao222_1 \U1811/U18/U1/U1  ( .x(net176), .a(net162), .b(pkt_done), .c(
        net162), .d(net176), .e(pkt_done), .f(net176) );
    aoi222_1 \U1664/U28/U30/U1  ( .x(\U1664/x[3] ), .a(\ncd[7] ), .b(\ncd[6] ), 
        .c(\ncd[7] ), .d(\U1664/U28/Z ), .e(\ncd[6] ), .f(\U1664/U28/Z ) );
    inv_1 \U1664/U28/U30/Uinv  ( .x(\U1664/U28/Z ), .a(\U1664/x[3] ) );
    aoi222_1 \U1664/U32/U30/U1  ( .x(\U1664/x[0] ), .a(\ncd[1] ), .b(\ncd[0] ), 
        .c(\ncd[1] ), .d(\U1664/U32/Z ), .e(\ncd[0] ), .f(\U1664/U32/Z ) );
    inv_1 \U1664/U32/U30/Uinv  ( .x(\U1664/U32/Z ), .a(\U1664/x[0] ) );
    aoi222_1 \U1664/U29/U30/U1  ( .x(\U1664/x[2] ), .a(\ncd[5] ), .b(\ncd[4] ), 
        .c(\ncd[5] ), .d(\U1664/U29/Z ), .e(\ncd[4] ), .f(\U1664/U29/Z ) );
    inv_1 \U1664/U29/U30/Uinv  ( .x(\U1664/U29/Z ), .a(\U1664/x[2] ) );
    aoi222_1 \U1664/U33/U30/U1  ( .x(\U1664/y[0] ), .a(\U1664/x[1] ), .b(
        \U1664/x[0] ), .c(\U1664/x[1] ), .d(\U1664/U33/Z ), .e(\U1664/x[0] ), 
        .f(\U1664/U33/Z ) );
    inv_1 \U1664/U33/U30/Uinv  ( .x(\U1664/U33/Z ), .a(\U1664/y[0] ) );
    aoi222_1 \U1664/U30/U30/U1  ( .x(\U1664/y[1] ), .a(\U1664/x[3] ), .b(
        \U1664/x[2] ), .c(\U1664/x[3] ), .d(\U1664/U30/Z ), .e(\U1664/x[2] ), 
        .f(\U1664/U30/Z ) );
    inv_1 \U1664/U30/U30/Uinv  ( .x(\U1664/U30/Z ), .a(\U1664/y[1] ) );
    aoi222_1 \U1664/U31/U30/U1  ( .x(\U1664/x[1] ), .a(\ncd[3] ), .b(\ncd[2] ), 
        .c(\ncd[3] ), .d(\U1664/U31/Z ), .e(\ncd[2] ), .f(\U1664/U31/Z ) );
    inv_1 \U1664/U31/U30/Uinv  ( .x(\U1664/U31/Z ), .a(\U1664/x[1] ) );
    aoi222_1 \U1664/U37/U30/U1  ( .x(pullcd), .a(\U1664/y[0] ), .b(
        \U1664/y[1] ), .c(\U1664/y[0] ), .d(\U1664/U37/Z ), .e(\U1664/y[1] ), 
        .f(\U1664/U37/Z ) );
    inv_1 \U1664/U37/U30/Uinv  ( .x(\U1664/U37/Z ), .a(pullcd) );
    nor3_1 \U1697/U21/Unr  ( .x(\U1697/U21/nr ), .a(rnw[0]), .b(pkt_normal), 
        .c(net149) );
    nand3_1 \U1697/U21/Und  ( .x(\U1697/U21/nd ), .a(rnw[0]), .b(pkt_normal), 
        .c(net149) );
    oa21_1 \U1697/U21/U1  ( .x(\U1697/U21/n2 ), .a(\U1697/U21/n2 ), .b(
        \U1697/U21/nr ), .c(\U1697/U21/nd ) );
    inv_1 \U1697/U21/U3  ( .x(write), .a(\U1697/U21/n2 ) );
    nor3_1 \U307/U21/Unr  ( .x(\U307/U21/nr ), .a(net149), .b(net150), .c(
        statusack) );
    nand3_1 \U307/U21/Und  ( .x(\U307/U21/nd ), .a(net149), .b(net150), .c(
        statusack) );
    oa21_1 \U307/U21/U1  ( .x(\U307/U21/n2 ), .a(\U307/U21/n2 ), .b(
        \U307/U21/nr ), .c(\U307/U21/nd ) );
    inv_1 \U307/U21/U3  ( .x(notify), .a(\U307/U21/n2 ) );
    nor3_1 \U1698/Unr  ( .x(\U1698/nr ), .a(rnw[1]), .b(pkt_normal), .c(net149
        ) );
    nand3_1 \U1698/Und  ( .x(\U1698/nd ), .a(rnw[1]), .b(pkt_normal), .c(
        net149) );
    oa21_1 \U1698/U1  ( .x(\U1698/n2 ), .a(\U1698/n2 ), .b(\U1698/nr ), .c(
        \U1698/nd ) );
    inv_2 \U1698/U3  ( .x(read), .a(\U1698/n2 ) );
    and2_1 \U1756/U1754/U8  ( .x(n17), .a(\opc_h[0] ), .b(pkt_normal) );
    and2_1 \U1756/U1755/U8  ( .x(n18), .a(\opc_l[0] ), .b(pkt_normal) );
    and2_1 \U1800/U1754/U8  ( .x(rnw[1]), .a(net0187), .b(pkt_normal) );
    and2_1 \U1800/U1755/U8  ( .x(rnw[0]), .a(net0208), .b(pkt_normal) );
    and2_1 \U1758/U1754/U8  ( .x(status[1]), .a(\opc_h[0] ), .b(net150) );
    and2_1 \U1758/U1755/U8  ( .x(status[0]), .a(\opc_l[0] ), .b(net150) );
    buf_2 \I6/U1653  ( .x(\I6/latch ), .a(net173) );
    nor2_1 \I6/U264/U5  ( .x(\I6/nlocalcd ), .a(reset), .b(\I6/localcd ) );
    nor2_1 \I6/U1659_0_/U5  ( .x(\I6/ncd[0] ), .a(\opc_l[0] ), .b(\opc_h[0] )
         );
    nor2_1 \I6/U1659_1_/U5  ( .x(\I6/ncd[1] ), .a(\opc_l[1] ), .b(\opc_h[1] )
         );
    nor2_1 \I6/U1659_2_/U5  ( .x(\I6/ncd[2] ), .a(\opc_l[2] ), .b(\I6/oh[2] )
         );
    nor2_1 \I6/U1659_3_/U5  ( .x(\I6/ncd[3] ), .a(\I6/ol[3] ), .b(\I6/oh[3] )
         );
    nor2_1 \I6/U1659_4_/U5  ( .x(\I6/ncd[4] ), .a(\I6/ol[4] ), .b(\I6/oh[4] )
         );
    nor2_1 \I6/U1659_5_/U5  ( .x(\I6/ncd[5] ), .a(net0208), .b(net0187) );
    nor2_1 \I6/U1659_6_/U5  ( .x(\I6/ncd[6] ), .a(\I6/ol[6] ), .b(\I6/oh[6] )
         );
    nor2_1 \I6/U1659_7_/U5  ( .x(\I6/ncd[7] ), .a(\I6/ol[7] ), .b(\I6/oh[7] )
         );
    nor2_1 \I6/U3/U5  ( .x(\I6/ctrlack_internal ), .a(\I6/acb ), .b(\I6/ba )
         );
    buf_2 \I6/U1665/U7  ( .x(\I6/driveh ), .a(net139) );
    buf_2 \I6/U1666/U7  ( .x(\I6/drivel ), .a(net139) );
    ao23_1 \I6/U1658_0_/U21/U1/U1  ( .x(\opc_l[0] ), .a(\I6/driveh ), .b(
        \opc_l[0] ), .c(\I6/driveh ), .d(cbl[0]), .e(n12) );
    ao23_1 \I6/U1658_1_/U21/U1/U1  ( .x(\opc_l[1] ), .a(\I6/driveh ), .b(
        \opc_l[1] ), .c(\I6/drivel ), .d(cbl[1]), .e(n12) );
    ao23_1 \I6/U1658_2_/U21/U1/U1  ( .x(\opc_l[2] ), .a(\I6/drivel ), .b(
        \opc_l[2] ), .c(n13), .d(cbl[2]), .e(n12) );
    ao23_1 \I6/U1658_3_/U21/U1/U1  ( .x(\I6/ol[3] ), .a(\I6/drivel ), .b(
        \I6/ol[3] ), .c(\I6/drivel ), .d(cbl[3]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_4_/U21/U1/U1  ( .x(\I6/ol[4] ), .a(n13), .b(\I6/ol[4] ), 
        .c(n13), .d(cbl[4]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_5_/U21/U1/U1  ( .x(net0208), .a(\I6/driveh ), .b(net0208), 
        .c(\I6/driveh ), .d(cbl[5]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_6_/U21/U1/U1  ( .x(\I6/ol[6] ), .a(n13), .b(\I6/ol[6] ), 
        .c(n13), .d(cbl[6]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_7_/U21/U1/U1  ( .x(\I6/ol[7] ), .a(n13), .b(\I6/ol[7] ), 
        .c(\I6/driveh ), .d(cbl[7]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_0_/U21/U1/U1  ( .x(\opc_h[0] ), .a(n13), .b(\opc_h[0] ), 
        .c(\I6/drivel ), .d(cbh[0]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_1_/U21/U1/U1  ( .x(\opc_h[1] ), .a(\I6/driveh ), .b(
        \opc_h[1] ), .c(n13), .d(cbh[1]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_2_/U21/U1/U1  ( .x(\I6/oh[2] ), .a(\I6/driveh ), .b(
        \I6/oh[2] ), .c(n13), .d(cbh[2]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_3_/U21/U1/U1  ( .x(\I6/oh[3] ), .a(\I6/drivel ), .b(
        \I6/oh[3] ), .c(\I6/drivel ), .d(cbh[3]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_4_/U21/U1/U1  ( .x(\I6/oh[4] ), .a(n13), .b(\I6/oh[4] ), 
        .c(\I6/driveh ), .d(cbh[4]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_5_/U21/U1/U1  ( .x(net0187), .a(\I6/driveh ), .b(net0187), 
        .c(\I6/driveh ), .d(cbh[5]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_6_/U21/U1/U1  ( .x(\I6/oh[6] ), .a(\I6/drivel ), .b(
        \I6/oh[6] ), .c(\I6/drivel ), .d(cbh[6]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_7_/U21/U1/U1  ( .x(\I6/oh[7] ), .a(\I6/drivel ), .b(
        \I6/oh[7] ), .c(n13), .d(cbh[7]), .e(\I6/latch ) );
    aoai211_1 \I6/U4/U28/U1/U1  ( .x(\I6/U4/U28/U1/clr ), .a(net139), .b(
        \I6/acb ), .c(\I6/nlocalcd ), .d(net173) );
    nand3_1 \I6/U4/U28/U1/U2  ( .x(\I6/U4/U28/U1/set ), .a(\I6/nlocalcd ), .b(
        net139), .c(\I6/acb ) );
    nand2_2 \I6/U4/U28/U1/U3  ( .x(net173), .a(\I6/U4/U28/U1/clr ), .b(
        \I6/U4/U28/U1/set ) );
    oai21_1 \I6/U1/U30/U1/U1  ( .x(\I6/acb ), .a(\I6/U1/Z ), .b(\I6/ba ), .c(
        net139) );
    inv_1 \I6/U1/U30/U1/U2  ( .x(\I6/U1/Z ), .a(\I6/acb ) );
    ao222_1 \I6/U5/U18/U1/U1  ( .x(\I6/ba ), .a(\I6/latch ), .b(n14), .c(
        \I6/latch ), .d(\I6/ba ), .e(n14), .f(\I6/ba ) );
    aoi222_1 \I6/U1664/U28/U30/U1  ( .x(\I6/U1664/x[3] ), .a(\I6/ncd[7] ), .b(
        \I6/ncd[6] ), .c(\I6/ncd[7] ), .d(\I6/U1664/U28/Z ), .e(\I6/ncd[6] ), 
        .f(\I6/U1664/U28/Z ) );
    inv_1 \I6/U1664/U28/U30/Uinv  ( .x(\I6/U1664/U28/Z ), .a(\I6/U1664/x[3] )
         );
    aoi222_1 \I6/U1664/U32/U30/U1  ( .x(\I6/U1664/x[0] ), .a(\I6/ncd[1] ), .b(
        \I6/ncd[0] ), .c(\I6/ncd[1] ), .d(\I6/U1664/U32/Z ), .e(\I6/ncd[0] ), 
        .f(\I6/U1664/U32/Z ) );
    inv_1 \I6/U1664/U32/U30/Uinv  ( .x(\I6/U1664/U32/Z ), .a(\I6/U1664/x[0] )
         );
    aoi222_1 \I6/U1664/U29/U30/U1  ( .x(\I6/U1664/x[2] ), .a(\I6/ncd[5] ), .b(
        \I6/ncd[4] ), .c(\I6/ncd[5] ), .d(\I6/U1664/U29/Z ), .e(\I6/ncd[4] ), 
        .f(\I6/U1664/U29/Z ) );
    inv_1 \I6/U1664/U29/U30/Uinv  ( .x(\I6/U1664/U29/Z ), .a(\I6/U1664/x[2] )
         );
    aoi222_1 \I6/U1664/U33/U30/U1  ( .x(\I6/U1664/y[0] ), .a(\I6/U1664/x[1] ), 
        .b(\I6/U1664/x[0] ), .c(\I6/U1664/x[1] ), .d(\I6/U1664/U33/Z ), .e(
        \I6/U1664/x[0] ), .f(\I6/U1664/U33/Z ) );
    inv_1 \I6/U1664/U33/U30/Uinv  ( .x(\I6/U1664/U33/Z ), .a(\I6/U1664/y[0] )
         );
    aoi222_1 \I6/U1664/U30/U30/U1  ( .x(\I6/U1664/y[1] ), .a(\I6/U1664/x[3] ), 
        .b(\I6/U1664/x[2] ), .c(\I6/U1664/x[3] ), .d(\I6/U1664/U30/Z ), .e(
        \I6/U1664/x[2] ), .f(\I6/U1664/U30/Z ) );
    inv_1 \I6/U1664/U30/U30/Uinv  ( .x(\I6/U1664/U30/Z ), .a(\I6/U1664/y[1] )
         );
    aoi222_1 \I6/U1664/U31/U30/U1  ( .x(\I6/U1664/x[1] ), .a(\I6/ncd[3] ), .b(
        \I6/ncd[2] ), .c(\I6/ncd[3] ), .d(\I6/U1664/U31/Z ), .e(\I6/ncd[2] ), 
        .f(\I6/U1664/U31/Z ) );
    inv_1 \I6/U1664/U31/U30/Uinv  ( .x(\I6/U1664/U31/Z ), .a(\I6/U1664/x[1] )
         );
    aoi222_1 \I6/U1664/U37/U30/U1  ( .x(\I6/localcd ), .a(\I6/U1664/y[0] ), 
        .b(\I6/U1664/y[1] ), .c(\I6/U1664/y[0] ), .d(\I6/U1664/U37/Z ), .e(
        \I6/U1664/y[1] ), .f(\I6/U1664/U37/Z ) );
    inv_1 \I6/U1664/U37/U30/Uinv  ( .x(\I6/U1664/U37/Z ), .a(\I6/localcd ) );
    nor3_1 \I6/U1669/Unr  ( .x(\I6/U1669/nr ), .a(\I6/ctrlack_internal ), .b(
        n13), .c(\I6/drivel ) );
    nand3_1 \I6/U1669/Und  ( .x(\I6/U1669/nd ), .a(\I6/ctrlack_internal ), .b(
        \I6/driveh ), .c(\I6/drivel ) );
    oa21_1 \I6/U1669/U1  ( .x(\I6/U1669/n2 ), .a(\I6/U1669/n2 ), .b(
        \I6/U1669/nr ), .c(\I6/U1669/nd ) );
    inv_2 \I6/U1669/U3  ( .x(net149), .a(\I6/U1669/n2 ) );
    buf_2 \U1667/U1653  ( .x(\U1667/latch ), .a(net167) );
    nor2_1 \U1667/U264/U5  ( .x(\U1667/nlocalcd ), .a(reset), .b(
        \U1667/localcd ) );
    nor2_1 \U1667/U1659_0_/U5  ( .x(\U1667/ncd[0] ), .a(rd[0]), .b(rd[32]) );
    nor2_1 \U1667/U1659_1_/U5  ( .x(\U1667/ncd[1] ), .a(rd[1]), .b(rd[33]) );
    nor2_1 \U1667/U1659_2_/U5  ( .x(\U1667/ncd[2] ), .a(rd[2]), .b(rd[34]) );
    nor2_1 \U1667/U1659_3_/U5  ( .x(\U1667/ncd[3] ), .a(rd[3]), .b(rd[35]) );
    nor2_1 \U1667/U1659_4_/U5  ( .x(\U1667/ncd[4] ), .a(rd[4]), .b(rd[36]) );
    nor2_1 \U1667/U1659_5_/U5  ( .x(\U1667/ncd[5] ), .a(rd[5]), .b(rd[37]) );
    nor2_1 \U1667/U1659_6_/U5  ( .x(\U1667/ncd[6] ), .a(rd[6]), .b(rd[38]) );
    nor2_1 \U1667/U1659_7_/U5  ( .x(\U1667/ncd[7] ), .a(rd[7]), .b(rd[39]) );
    nor2_1 \U1667/U3/U5  ( .x(\U1667/ctrlack_internal ), .a(\U1667/acb ), .b(
        \U1667/ba ) );
    buf_2 \U1667/U1665/U7  ( .x(\U1667/driveh ), .a(read_lhw) );
    buf_2 \U1667/U1666/U7  ( .x(\U1667/drivel ), .a(read_lhw) );
    ao23_1 \U1667/U1658_0_/U21/U1/U1  ( .x(rd[0]), .a(n11), .b(rd[0]), .c(
        \U1667/drivel ), .d(cbl[0]), .e(n10) );
    ao23_1 \U1667/U1658_1_/U21/U1/U1  ( .x(rd[1]), .a(n11), .b(rd[1]), .c(
        \U1667/driveh ), .d(cbl[1]), .e(n10) );
    ao23_1 \U1667/U1658_2_/U21/U1/U1  ( .x(rd[2]), .a(\U1667/driveh ), .b(rd
        [2]), .c(n11), .d(cbl[2]), .e(n10) );
    ao23_1 \U1667/U1658_3_/U21/U1/U1  ( .x(rd[3]), .a(n11), .b(rd[3]), .c(
        \U1667/driveh ), .d(cbl[3]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_4_/U21/U1/U1  ( .x(rd[4]), .a(\U1667/drivel ), .b(rd
        [4]), .c(n11), .d(cbl[4]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_5_/U21/U1/U1  ( .x(rd[5]), .a(\U1667/drivel ), .b(rd
        [5]), .c(n11), .d(cbl[5]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_6_/U21/U1/U1  ( .x(rd[6]), .a(\U1667/driveh ), .b(rd
        [6]), .c(\U1667/drivel ), .d(cbl[6]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_7_/U21/U1/U1  ( .x(rd[7]), .a(\U1667/driveh ), .b(rd
        [7]), .c(\U1667/driveh ), .d(cbl[7]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_0_/U21/U1/U1  ( .x(rd[32]), .a(\U1667/drivel ), .b(rd
        [32]), .c(n11), .d(cbh[0]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_1_/U21/U1/U1  ( .x(rd[33]), .a(\U1667/driveh ), .b(rd
        [33]), .c(\U1667/drivel ), .d(cbh[1]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_2_/U21/U1/U1  ( .x(rd[34]), .a(\U1667/drivel ), .b(rd
        [34]), .c(\U1667/drivel ), .d(cbh[2]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_3_/U21/U1/U1  ( .x(rd[35]), .a(\U1667/driveh ), .b(rd
        [35]), .c(\U1667/driveh ), .d(cbh[3]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_4_/U21/U1/U1  ( .x(rd[36]), .a(\U1667/drivel ), .b(rd
        [36]), .c(\U1667/driveh ), .d(cbh[4]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_5_/U21/U1/U1  ( .x(rd[37]), .a(\U1667/driveh ), .b(rd
        [37]), .c(n11), .d(cbh[5]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_6_/U21/U1/U1  ( .x(rd[38]), .a(n11), .b(rd[38]), .c(
        \U1667/drivel ), .d(cbh[6]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_7_/U21/U1/U1  ( .x(rd[39]), .a(n11), .b(rd[39]), .c(
        n11), .d(cbh[7]), .e(\U1667/latch ) );
    aoai211_1 \U1667/U4/U28/U1/U1  ( .x(\U1667/U4/U28/U1/clr ), .a(read_lhw), 
        .b(\U1667/acb ), .c(\U1667/nlocalcd ), .d(net167) );
    nand3_1 \U1667/U4/U28/U1/U2  ( .x(\U1667/U4/U28/U1/set ), .a(
        \U1667/nlocalcd ), .b(read_lhw), .c(\U1667/acb ) );
    nand2_2 \U1667/U4/U28/U1/U3  ( .x(net167), .a(\U1667/U4/U28/U1/clr ), .b(
        \U1667/U4/U28/U1/set ) );
    oai21_1 \U1667/U1/U30/U1/U1  ( .x(\U1667/acb ), .a(\U1667/U1/Z ), .b(
        \U1667/ba ), .c(read_lhw) );
    inv_1 \U1667/U1/U30/U1/U2  ( .x(\U1667/U1/Z ), .a(\U1667/acb ) );
    ao222_1 \U1667/U5/U18/U1/U1  ( .x(\U1667/ba ), .a(\U1667/latch ), .b(n14), 
        .c(\U1667/latch ), .d(\U1667/ba ), .e(n14), .f(\U1667/ba ) );
    aoi222_1 \U1667/U1664/U28/U30/U1  ( .x(\U1667/U1664/x[3] ), .a(
        \U1667/ncd[7] ), .b(\U1667/ncd[6] ), .c(\U1667/ncd[7] ), .d(
        \U1667/U1664/U28/Z ), .e(\U1667/ncd[6] ), .f(\U1667/U1664/U28/Z ) );
    inv_1 \U1667/U1664/U28/U30/Uinv  ( .x(\U1667/U1664/U28/Z ), .a(
        \U1667/U1664/x[3] ) );
    aoi222_1 \U1667/U1664/U32/U30/U1  ( .x(\U1667/U1664/x[0] ), .a(
        \U1667/ncd[1] ), .b(\U1667/ncd[0] ), .c(\U1667/ncd[1] ), .d(
        \U1667/U1664/U32/Z ), .e(\U1667/ncd[0] ), .f(\U1667/U1664/U32/Z ) );
    inv_1 \U1667/U1664/U32/U30/Uinv  ( .x(\U1667/U1664/U32/Z ), .a(
        \U1667/U1664/x[0] ) );
    aoi222_1 \U1667/U1664/U29/U30/U1  ( .x(\U1667/U1664/x[2] ), .a(
        \U1667/ncd[5] ), .b(\U1667/ncd[4] ), .c(\U1667/ncd[5] ), .d(
        \U1667/U1664/U29/Z ), .e(\U1667/ncd[4] ), .f(\U1667/U1664/U29/Z ) );
    inv_1 \U1667/U1664/U29/U30/Uinv  ( .x(\U1667/U1664/U29/Z ), .a(
        \U1667/U1664/x[2] ) );
    aoi222_1 \U1667/U1664/U33/U30/U1  ( .x(\U1667/U1664/y[0] ), .a(
        \U1667/U1664/x[1] ), .b(\U1667/U1664/x[0] ), .c(\U1667/U1664/x[1] ), 
        .d(\U1667/U1664/U33/Z ), .e(\U1667/U1664/x[0] ), .f(
        \U1667/U1664/U33/Z ) );
    inv_1 \U1667/U1664/U33/U30/Uinv  ( .x(\U1667/U1664/U33/Z ), .a(
        \U1667/U1664/y[0] ) );
    aoi222_1 \U1667/U1664/U30/U30/U1  ( .x(\U1667/U1664/y[1] ), .a(
        \U1667/U1664/x[3] ), .b(\U1667/U1664/x[2] ), .c(\U1667/U1664/x[3] ), 
        .d(\U1667/U1664/U30/Z ), .e(\U1667/U1664/x[2] ), .f(
        \U1667/U1664/U30/Z ) );
    inv_1 \U1667/U1664/U30/U30/Uinv  ( .x(\U1667/U1664/U30/Z ), .a(
        \U1667/U1664/y[1] ) );
    aoi222_1 \U1667/U1664/U31/U30/U1  ( .x(\U1667/U1664/x[1] ), .a(
        \U1667/ncd[3] ), .b(\U1667/ncd[2] ), .c(\U1667/ncd[3] ), .d(
        \U1667/U1664/U31/Z ), .e(\U1667/ncd[2] ), .f(\U1667/U1664/U31/Z ) );
    inv_1 \U1667/U1664/U31/U30/Uinv  ( .x(\U1667/U1664/U31/Z ), .a(
        \U1667/U1664/x[1] ) );
    aoi222_1 \U1667/U1664/U37/U30/U1  ( .x(\U1667/localcd ), .a(
        \U1667/U1664/y[0] ), .b(\U1667/U1664/y[1] ), .c(\U1667/U1664/y[0] ), 
        .d(\U1667/U1664/U37/Z ), .e(\U1667/U1664/y[1] ), .f(
        \U1667/U1664/U37/Z ) );
    inv_1 \U1667/U1664/U37/U30/Uinv  ( .x(\U1667/U1664/U37/Z ), .a(
        \U1667/localcd ) );
    nor3_1 \U1667/U1669/Unr  ( .x(\U1667/U1669/nr ), .a(
        \U1667/ctrlack_internal ), .b(n11), .c(\U1667/drivel ) );
    nand3_1 \U1667/U1669/Und  ( .x(\U1667/U1669/nd ), .a(
        \U1667/ctrlack_internal ), .b(\U1667/driveh ), .c(\U1667/drivel ) );
    oa21_1 \U1667/U1669/U1  ( .x(\U1667/U1669/n2 ), .a(\U1667/U1669/n2 ), .b(
        \U1667/U1669/nr ), .c(\U1667/U1669/nd ) );
    inv_2 \U1667/U1669/U3  ( .x(net193), .a(\U1667/U1669/n2 ) );
    buf_2 \U1650/U1653  ( .x(\U1650/latch ), .a(net172) );
    nor2_1 \U1650/U264/U5  ( .x(\U1650/nlocalcd ), .a(reset), .b(
        \U1650/localcd ) );
    nor2_1 \U1650/U1659_0_/U5  ( .x(\U1650/ncd[0] ), .a(\U1650/ol[0] ), .b(
        \U1650/oh[0] ) );
    nor2_1 \U1650/U1659_1_/U5  ( .x(\U1650/ncd[1] ), .a(\U1650/ol[1] ), .b(
        \U1650/oh[1] ) );
    nor2_1 \U1650/U1659_2_/U5  ( .x(\U1650/ncd[2] ), .a(\U1650/ol[2] ), .b(
        \U1650/oh[2] ) );
    nor2_1 \U1650/U1659_3_/U5  ( .x(\U1650/ncd[3] ), .a(\U1650/ol[3] ), .b(
        \U1650/oh[3] ) );
    nor2_1 \U1650/U1659_4_/U5  ( .x(\U1650/ncd[4] ), .a(\U1650/ol[4] ), .b(
        \U1650/oh[4] ) );
    nor2_1 \U1650/U1659_5_/U5  ( .x(\U1650/ncd[5] ), .a(\col_l[0] ), .b(
        \col_h[0] ) );
    nor2_1 \U1650/U1659_6_/U5  ( .x(\U1650/ncd[6] ), .a(\col_l[1] ), .b(
        \col_h[1] ) );
    nor2_1 \U1650/U1659_7_/U5  ( .x(\U1650/ncd[7] ), .a(\col_l[2] ), .b(
        \col_h[2] ) );
    nor2_1 \U1650/U3/U5  ( .x(\U1650/ctrlack_internal ), .a(\U1650/acb ), .b(
        \U1650/ba ) );
    buf_2 \U1650/U1665/U7  ( .x(\U1650/driveh ), .a(start_receiving) );
    buf_2 \U1650/U1666/U7  ( .x(\U1650/drivel ), .a(start_receiving) );
    ao23_1 \U1650/U1658_0_/U21/U1/U1  ( .x(\U1650/ol[0] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[0] ), .c(\U1650/drivel ), .d(cbl[0]), .e(n7) );
    ao23_1 \U1650/U1658_1_/U21/U1/U1  ( .x(\U1650/ol[1] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[1] ), .c(\U1650/drivel ), .d(cbl[1]), .e(n7) );
    ao23_1 \U1650/U1658_2_/U21/U1/U1  ( .x(\U1650/ol[2] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[2] ), .c(\U1650/drivel ), .d(cbl[2]), .e(n7) );
    ao23_1 \U1650/U1658_3_/U21/U1/U1  ( .x(\U1650/ol[3] ), .a(n9), .b(
        \U1650/ol[3] ), .c(\U1650/drivel ), .d(cbl[3]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1658_4_/U21/U1/U1  ( .x(\U1650/ol[4] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[4] ), .c(\U1650/drivel ), .d(cbl[4]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1658_5_/U21/U1/U1  ( .x(\col_l[0] ), .a(\U1650/drivel ), 
        .b(\col_l[0] ), .c(\U1650/drivel ), .d(cbl[5]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1658_6_/U21/U1/U1  ( .x(\col_l[1] ), .a(n9), .b(\col_l[1] ), 
        .c(\U1650/drivel ), .d(cbl[6]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1658_7_/U21/U1/U1  ( .x(\col_l[2] ), .a(n9), .b(\col_l[2] ), 
        .c(\U1650/drivel ), .d(cbl[7]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_0_/U21/U1/U1  ( .x(\U1650/oh[0] ), .a(\U1650/driveh ), 
        .b(\U1650/oh[0] ), .c(\U1650/driveh ), .d(cbh[0]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1651_1_/U21/U1/U1  ( .x(\U1650/oh[1] ), .a(\U1650/driveh ), 
        .b(\U1650/oh[1] ), .c(\U1650/driveh ), .d(cbh[1]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1651_2_/U21/U1/U1  ( .x(\U1650/oh[2] ), .a(\U1650/driveh ), 
        .b(\U1650/oh[2] ), .c(\U1650/driveh ), .d(cbh[2]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1651_3_/U21/U1/U1  ( .x(\U1650/oh[3] ), .a(n8), .b(
        \U1650/oh[3] ), .c(\U1650/driveh ), .d(cbh[3]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_4_/U21/U1/U1  ( .x(\U1650/oh[4] ), .a(n8), .b(
        \U1650/oh[4] ), .c(\U1650/driveh ), .d(cbh[4]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_5_/U21/U1/U1  ( .x(\col_h[0] ), .a(\U1650/driveh ), 
        .b(\col_h[0] ), .c(\U1650/driveh ), .d(cbh[5]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_6_/U21/U1/U1  ( .x(\col_h[1] ), .a(n8), .b(\col_h[1] ), 
        .c(\U1650/driveh ), .d(cbh[6]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_7_/U21/U1/U1  ( .x(\col_h[2] ), .a(\U1650/driveh ), 
        .b(\col_h[2] ), .c(\U1650/driveh ), .d(cbh[7]), .e(\U1650/latch ) );
    aoai211_1 \U1650/U4/U28/U1/U1  ( .x(\U1650/U4/U28/U1/clr ), .a(
        start_receiving), .b(\U1650/acb ), .c(\U1650/nlocalcd ), .d(net172) );
    nand3_1 \U1650/U4/U28/U1/U2  ( .x(\U1650/U4/U28/U1/set ), .a(
        \U1650/nlocalcd ), .b(start_receiving), .c(\U1650/acb ) );
    nand2_2 \U1650/U4/U28/U1/U3  ( .x(net172), .a(\U1650/U4/U28/U1/clr ), .b(
        \U1650/U4/U28/U1/set ) );
    oai21_1 \U1650/U1/U30/U1/U1  ( .x(\U1650/acb ), .a(\U1650/U1/Z ), .b(
        \U1650/ba ), .c(start_receiving) );
    inv_1 \U1650/U1/U30/U1/U2  ( .x(\U1650/U1/Z ), .a(\U1650/acb ) );
    ao222_1 \U1650/U5/U18/U1/U1  ( .x(\U1650/ba ), .a(\U1650/latch ), .b(n14), 
        .c(\U1650/latch ), .d(\U1650/ba ), .e(n14), .f(\U1650/ba ) );
    aoi222_1 \U1650/U1664/U28/U30/U1  ( .x(\U1650/U1664/x[3] ), .a(
        \U1650/ncd[7] ), .b(\U1650/ncd[6] ), .c(\U1650/ncd[7] ), .d(
        \U1650/U1664/U28/Z ), .e(\U1650/ncd[6] ), .f(\U1650/U1664/U28/Z ) );
    inv_1 \U1650/U1664/U28/U30/Uinv  ( .x(\U1650/U1664/U28/Z ), .a(
        \U1650/U1664/x[3] ) );
    aoi222_1 \U1650/U1664/U32/U30/U1  ( .x(\U1650/U1664/x[0] ), .a(
        \U1650/ncd[1] ), .b(\U1650/ncd[0] ), .c(\U1650/ncd[1] ), .d(
        \U1650/U1664/U32/Z ), .e(\U1650/ncd[0] ), .f(\U1650/U1664/U32/Z ) );
    inv_1 \U1650/U1664/U32/U30/Uinv  ( .x(\U1650/U1664/U32/Z ), .a(
        \U1650/U1664/x[0] ) );
    aoi222_1 \U1650/U1664/U29/U30/U1  ( .x(\U1650/U1664/x[2] ), .a(
        \U1650/ncd[5] ), .b(\U1650/ncd[4] ), .c(\U1650/ncd[5] ), .d(
        \U1650/U1664/U29/Z ), .e(\U1650/ncd[4] ), .f(\U1650/U1664/U29/Z ) );
    inv_1 \U1650/U1664/U29/U30/Uinv  ( .x(\U1650/U1664/U29/Z ), .a(
        \U1650/U1664/x[2] ) );
    aoi222_1 \U1650/U1664/U33/U30/U1  ( .x(\U1650/U1664/y[0] ), .a(
        \U1650/U1664/x[1] ), .b(\U1650/U1664/x[0] ), .c(\U1650/U1664/x[1] ), 
        .d(\U1650/U1664/U33/Z ), .e(\U1650/U1664/x[0] ), .f(
        \U1650/U1664/U33/Z ) );
    inv_1 \U1650/U1664/U33/U30/Uinv  ( .x(\U1650/U1664/U33/Z ), .a(
        \U1650/U1664/y[0] ) );
    aoi222_1 \U1650/U1664/U30/U30/U1  ( .x(\U1650/U1664/y[1] ), .a(
        \U1650/U1664/x[3] ), .b(\U1650/U1664/x[2] ), .c(\U1650/U1664/x[3] ), 
        .d(\U1650/U1664/U30/Z ), .e(\U1650/U1664/x[2] ), .f(
        \U1650/U1664/U30/Z ) );
    inv_1 \U1650/U1664/U30/U30/Uinv  ( .x(\U1650/U1664/U30/Z ), .a(
        \U1650/U1664/y[1] ) );
    aoi222_1 \U1650/U1664/U31/U30/U1  ( .x(\U1650/U1664/x[1] ), .a(
        \U1650/ncd[3] ), .b(\U1650/ncd[2] ), .c(\U1650/ncd[3] ), .d(
        \U1650/U1664/U31/Z ), .e(\U1650/ncd[2] ), .f(\U1650/U1664/U31/Z ) );
    inv_1 \U1650/U1664/U31/U30/Uinv  ( .x(\U1650/U1664/U31/Z ), .a(
        \U1650/U1664/x[1] ) );
    aoi222_1 \U1650/U1664/U37/U30/U1  ( .x(\U1650/localcd ), .a(
        \U1650/U1664/y[0] ), .b(\U1650/U1664/y[1] ), .c(\U1650/U1664/y[0] ), 
        .d(\U1650/U1664/U37/Z ), .e(\U1650/U1664/y[1] ), .f(
        \U1650/U1664/U37/Z ) );
    inv_1 \U1650/U1664/U37/U30/Uinv  ( .x(\U1650/U1664/U37/Z ), .a(
        \U1650/localcd ) );
    nor3_1 \U1650/U1669/Unr  ( .x(\U1650/U1669/nr ), .a(
        \U1650/ctrlack_internal ), .b(\U1650/drivel ), .c(\U1650/driveh ) );
    nand3_1 \U1650/U1669/Und  ( .x(\U1650/U1669/nd ), .a(
        \U1650/ctrlack_internal ), .b(\U1650/drivel ), .c(\U1650/driveh ) );
    oa21_1 \U1650/U1669/U1  ( .x(\U1650/U1669/n2 ), .a(\U1650/U1669/n2 ), .b(
        \U1650/U1669/nr ), .c(\U1650/U1669/nd ) );
    inv_2 \U1650/U1669/U3  ( .x(net139), .a(\U1650/U1669/n2 ) );
    buf_2 \U1666/U1653  ( .x(\U1666/latch ), .a(net169) );
    nor2_1 \U1666/U264/U5  ( .x(\U1666/nlocalcd ), .a(reset), .b(
        \U1666/localcd ) );
    nor2_1 \U1666/U1659_0_/U5  ( .x(\U1666/ncd[0] ), .a(rd[24]), .b(rd[56]) );
    nor2_1 \U1666/U1659_1_/U5  ( .x(\U1666/ncd[1] ), .a(rd[25]), .b(rd[57]) );
    nor2_1 \U1666/U1659_2_/U5  ( .x(\U1666/ncd[2] ), .a(rd[26]), .b(rd[58]) );
    nor2_1 \U1666/U1659_3_/U5  ( .x(\U1666/ncd[3] ), .a(rd[27]), .b(rd[59]) );
    nor2_1 \U1666/U1659_4_/U5  ( .x(\U1666/ncd[4] ), .a(rd[28]), .b(rd[60]) );
    nor2_1 \U1666/U1659_5_/U5  ( .x(\U1666/ncd[5] ), .a(rd[29]), .b(rd[61]) );
    nor2_1 \U1666/U1659_6_/U5  ( .x(\U1666/ncd[6] ), .a(rd[30]), .b(rd[62]) );
    nor2_1 \U1666/U1659_7_/U5  ( .x(\U1666/ncd[7] ), .a(rd[31]), .b(rd[63]) );
    nor2_1 \U1666/U3/U5  ( .x(\U1666/ctrlack_internal ), .a(\U1666/acb ), .b(
        \U1666/ba ) );
    buf_2 \U1666/U1665/U7  ( .x(\U1666/driveh ), .a(read) );
    buf_2 \U1666/U1666/U7  ( .x(\U1666/drivel ), .a(read) );
    ao23_1 \U1666/U1658_0_/U21/U1/U1  ( .x(rd[24]), .a(n6), .b(rd[24]), .c(
        \U1666/drivel ), .d(cbl[0]), .e(n5) );
    ao23_1 \U1666/U1658_1_/U21/U1/U1  ( .x(rd[25]), .a(n6), .b(rd[25]), .c(
        \U1666/driveh ), .d(cbl[1]), .e(n5) );
    ao23_1 \U1666/U1658_2_/U21/U1/U1  ( .x(rd[26]), .a(\U1666/driveh ), .b(rd
        [26]), .c(n6), .d(cbl[2]), .e(n5) );
    ao23_1 \U1666/U1658_3_/U21/U1/U1  ( .x(rd[27]), .a(n6), .b(rd[27]), .c(
        \U1666/driveh ), .d(cbl[3]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_4_/U21/U1/U1  ( .x(rd[28]), .a(\U1666/drivel ), .b(rd
        [28]), .c(n6), .d(cbl[4]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_5_/U21/U1/U1  ( .x(rd[29]), .a(\U1666/drivel ), .b(rd
        [29]), .c(n6), .d(cbl[5]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_6_/U21/U1/U1  ( .x(rd[30]), .a(\U1666/driveh ), .b(rd
        [30]), .c(\U1666/drivel ), .d(cbl[6]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_7_/U21/U1/U1  ( .x(rd[31]), .a(\U1666/driveh ), .b(rd
        [31]), .c(\U1666/driveh ), .d(cbl[7]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_0_/U21/U1/U1  ( .x(rd[56]), .a(\U1666/drivel ), .b(rd
        [56]), .c(n6), .d(cbh[0]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_1_/U21/U1/U1  ( .x(rd[57]), .a(\U1666/driveh ), .b(rd
        [57]), .c(\U1666/drivel ), .d(cbh[1]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_2_/U21/U1/U1  ( .x(rd[58]), .a(\U1666/drivel ), .b(rd
        [58]), .c(\U1666/drivel ), .d(cbh[2]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_3_/U21/U1/U1  ( .x(rd[59]), .a(\U1666/driveh ), .b(rd
        [59]), .c(\U1666/driveh ), .d(cbh[3]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_4_/U21/U1/U1  ( .x(rd[60]), .a(\U1666/drivel ), .b(rd
        [60]), .c(\U1666/driveh ), .d(cbh[4]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_5_/U21/U1/U1  ( .x(rd[61]), .a(\U1666/driveh ), .b(rd
        [61]), .c(n6), .d(cbh[5]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_6_/U21/U1/U1  ( .x(rd[62]), .a(n6), .b(rd[62]), .c(
        \U1666/drivel ), .d(cbh[6]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_7_/U21/U1/U1  ( .x(rd[63]), .a(n6), .b(rd[63]), .c(n6), 
        .d(cbh[7]), .e(\U1666/latch ) );
    aoai211_1 \U1666/U4/U28/U1/U1  ( .x(\U1666/U4/U28/U1/clr ), .a(read), .b(
        \U1666/acb ), .c(\U1666/nlocalcd ), .d(net169) );
    nand3_1 \U1666/U4/U28/U1/U2  ( .x(\U1666/U4/U28/U1/set ), .a(
        \U1666/nlocalcd ), .b(read), .c(\U1666/acb ) );
    nand2_2 \U1666/U4/U28/U1/U3  ( .x(net169), .a(\U1666/U4/U28/U1/clr ), .b(
        \U1666/U4/U28/U1/set ) );
    oai21_1 \U1666/U1/U30/U1/U1  ( .x(\U1666/acb ), .a(\U1666/U1/Z ), .b(
        \U1666/ba ), .c(read) );
    inv_1 \U1666/U1/U30/U1/U2  ( .x(\U1666/U1/Z ), .a(\U1666/acb ) );
    ao222_1 \U1666/U5/U18/U1/U1  ( .x(\U1666/ba ), .a(\U1666/latch ), .b(n14), 
        .c(\U1666/latch ), .d(\U1666/ba ), .e(n14), .f(\U1666/ba ) );
    aoi222_1 \U1666/U1664/U28/U30/U1  ( .x(\U1666/U1664/x[3] ), .a(
        \U1666/ncd[7] ), .b(\U1666/ncd[6] ), .c(\U1666/ncd[7] ), .d(
        \U1666/U1664/U28/Z ), .e(\U1666/ncd[6] ), .f(\U1666/U1664/U28/Z ) );
    inv_1 \U1666/U1664/U28/U30/Uinv  ( .x(\U1666/U1664/U28/Z ), .a(
        \U1666/U1664/x[3] ) );
    aoi222_1 \U1666/U1664/U32/U30/U1  ( .x(\U1666/U1664/x[0] ), .a(
        \U1666/ncd[1] ), .b(\U1666/ncd[0] ), .c(\U1666/ncd[1] ), .d(
        \U1666/U1664/U32/Z ), .e(\U1666/ncd[0] ), .f(\U1666/U1664/U32/Z ) );
    inv_1 \U1666/U1664/U32/U30/Uinv  ( .x(\U1666/U1664/U32/Z ), .a(
        \U1666/U1664/x[0] ) );
    aoi222_1 \U1666/U1664/U29/U30/U1  ( .x(\U1666/U1664/x[2] ), .a(
        \U1666/ncd[5] ), .b(\U1666/ncd[4] ), .c(\U1666/ncd[5] ), .d(
        \U1666/U1664/U29/Z ), .e(\U1666/ncd[4] ), .f(\U1666/U1664/U29/Z ) );
    inv_1 \U1666/U1664/U29/U30/Uinv  ( .x(\U1666/U1664/U29/Z ), .a(
        \U1666/U1664/x[2] ) );
    aoi222_1 \U1666/U1664/U33/U30/U1  ( .x(\U1666/U1664/y[0] ), .a(
        \U1666/U1664/x[1] ), .b(\U1666/U1664/x[0] ), .c(\U1666/U1664/x[1] ), 
        .d(\U1666/U1664/U33/Z ), .e(\U1666/U1664/x[0] ), .f(
        \U1666/U1664/U33/Z ) );
    inv_1 \U1666/U1664/U33/U30/Uinv  ( .x(\U1666/U1664/U33/Z ), .a(
        \U1666/U1664/y[0] ) );
    aoi222_1 \U1666/U1664/U30/U30/U1  ( .x(\U1666/U1664/y[1] ), .a(
        \U1666/U1664/x[3] ), .b(\U1666/U1664/x[2] ), .c(\U1666/U1664/x[3] ), 
        .d(\U1666/U1664/U30/Z ), .e(\U1666/U1664/x[2] ), .f(
        \U1666/U1664/U30/Z ) );
    inv_1 \U1666/U1664/U30/U30/Uinv  ( .x(\U1666/U1664/U30/Z ), .a(
        \U1666/U1664/y[1] ) );
    aoi222_1 \U1666/U1664/U31/U30/U1  ( .x(\U1666/U1664/x[1] ), .a(
        \U1666/ncd[3] ), .b(\U1666/ncd[2] ), .c(\U1666/ncd[3] ), .d(
        \U1666/U1664/U31/Z ), .e(\U1666/ncd[2] ), .f(\U1666/U1664/U31/Z ) );
    inv_1 \U1666/U1664/U31/U30/Uinv  ( .x(\U1666/U1664/U31/Z ), .a(
        \U1666/U1664/x[1] ) );
    aoi222_1 \U1666/U1664/U37/U30/U1  ( .x(\U1666/localcd ), .a(
        \U1666/U1664/y[0] ), .b(\U1666/U1664/y[1] ), .c(\U1666/U1664/y[0] ), 
        .d(\U1666/U1664/U37/Z ), .e(\U1666/U1664/y[1] ), .f(
        \U1666/U1664/U37/Z ) );
    inv_1 \U1666/U1664/U37/U30/Uinv  ( .x(\U1666/U1664/U37/Z ), .a(
        \U1666/localcd ) );
    nor3_1 \U1666/U1669/Unr  ( .x(\U1666/U1669/nr ), .a(
        \U1666/ctrlack_internal ), .b(n6), .c(\U1666/drivel ) );
    nand3_1 \U1666/U1669/Und  ( .x(\U1666/U1669/nd ), .a(
        \U1666/ctrlack_internal ), .b(\U1666/driveh ), .c(\U1666/drivel ) );
    oa21_1 \U1666/U1669/U1  ( .x(\U1666/U1669/n2 ), .a(\U1666/U1669/n2 ), .b(
        \U1666/U1669/nr ), .c(\U1666/U1669/nd ) );
    inv_2 \U1666/U1669/U3  ( .x(net94), .a(\U1666/U1669/n2 ) );
    buf_2 \I1/U1653  ( .x(\I1/latch ), .a(net166) );
    nor2_1 \I1/U264/U5  ( .x(\I1/nlocalcd ), .a(reset), .b(\I1/localcd ) );
    nor2_1 \I1/U1659_0_/U5  ( .x(\I1/ncd[0] ), .a(rd[8]), .b(rd[40]) );
    nor2_1 \I1/U1659_1_/U5  ( .x(\I1/ncd[1] ), .a(rd[9]), .b(rd[41]) );
    nor2_1 \I1/U1659_2_/U5  ( .x(\I1/ncd[2] ), .a(rd[10]), .b(rd[42]) );
    nor2_1 \I1/U1659_3_/U5  ( .x(\I1/ncd[3] ), .a(rd[11]), .b(rd[43]) );
    nor2_1 \I1/U1659_4_/U5  ( .x(\I1/ncd[4] ), .a(rd[12]), .b(rd[44]) );
    nor2_1 \I1/U1659_5_/U5  ( .x(\I1/ncd[5] ), .a(rd[13]), .b(rd[45]) );
    nor2_1 \I1/U1659_6_/U5  ( .x(\I1/ncd[6] ), .a(rd[14]), .b(rd[46]) );
    nor2_1 \I1/U1659_7_/U5  ( .x(\I1/ncd[7] ), .a(rd[15]), .b(rd[47]) );
    nor2_1 \I1/U3/U5  ( .x(\I1/ctrlack_internal ), .a(\I1/acb ), .b(\I1/ba )
         );
    buf_2 \I1/U1665/U7  ( .x(\I1/driveh ), .a(net103) );
    buf_2 \I1/U1666/U7  ( .x(\I1/drivel ), .a(net103) );
    ao23_1 \I1/U1658_0_/U21/U1/U1  ( .x(rd[8]), .a(n4), .b(rd[8]), .c(
        \I1/drivel ), .d(cbl[0]), .e(n3) );
    ao23_1 \I1/U1658_1_/U21/U1/U1  ( .x(rd[9]), .a(n4), .b(rd[9]), .c(
        \I1/driveh ), .d(cbl[1]), .e(n3) );
    ao23_1 \I1/U1658_2_/U21/U1/U1  ( .x(rd[10]), .a(\I1/driveh ), .b(rd[10]), 
        .c(n4), .d(cbl[2]), .e(n3) );
    ao23_1 \I1/U1658_3_/U21/U1/U1  ( .x(rd[11]), .a(n4), .b(rd[11]), .c(
        \I1/driveh ), .d(cbl[3]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_4_/U21/U1/U1  ( .x(rd[12]), .a(\I1/drivel ), .b(rd[12]), 
        .c(n4), .d(cbl[4]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_5_/U21/U1/U1  ( .x(rd[13]), .a(\I1/drivel ), .b(rd[13]), 
        .c(n4), .d(cbl[5]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_6_/U21/U1/U1  ( .x(rd[14]), .a(\I1/driveh ), .b(rd[14]), 
        .c(\I1/drivel ), .d(cbl[6]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_7_/U21/U1/U1  ( .x(rd[15]), .a(\I1/driveh ), .b(rd[15]), 
        .c(\I1/driveh ), .d(cbl[7]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_0_/U21/U1/U1  ( .x(rd[40]), .a(\I1/drivel ), .b(rd[40]), 
        .c(n4), .d(cbh[0]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_1_/U21/U1/U1  ( .x(rd[41]), .a(\I1/driveh ), .b(rd[41]), 
        .c(\I1/drivel ), .d(cbh[1]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_2_/U21/U1/U1  ( .x(rd[42]), .a(\I1/drivel ), .b(rd[42]), 
        .c(\I1/drivel ), .d(cbh[2]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_3_/U21/U1/U1  ( .x(rd[43]), .a(\I1/driveh ), .b(rd[43]), 
        .c(\I1/driveh ), .d(cbh[3]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_4_/U21/U1/U1  ( .x(rd[44]), .a(\I1/drivel ), .b(rd[44]), 
        .c(\I1/driveh ), .d(cbh[4]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_5_/U21/U1/U1  ( .x(rd[45]), .a(\I1/driveh ), .b(rd[45]), 
        .c(n4), .d(cbh[5]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_6_/U21/U1/U1  ( .x(rd[46]), .a(n4), .b(rd[46]), .c(
        \I1/drivel ), .d(cbh[6]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_7_/U21/U1/U1  ( .x(rd[47]), .a(n4), .b(rd[47]), .c(n4), 
        .d(cbh[7]), .e(\I1/latch ) );
    aoai211_1 \I1/U4/U28/U1/U1  ( .x(\I1/U4/U28/U1/clr ), .a(net103), .b(
        \I1/acb ), .c(\I1/nlocalcd ), .d(net166) );
    nand3_1 \I1/U4/U28/U1/U2  ( .x(\I1/U4/U28/U1/set ), .a(\I1/nlocalcd ), .b(
        net103), .c(\I1/acb ) );
    nand2_2 \I1/U4/U28/U1/U3  ( .x(net166), .a(\I1/U4/U28/U1/clr ), .b(
        \I1/U4/U28/U1/set ) );
    oai21_1 \I1/U1/U30/U1/U1  ( .x(\I1/acb ), .a(\I1/U1/Z ), .b(\I1/ba ), .c(
        net103) );
    inv_1 \I1/U1/U30/U1/U2  ( .x(\I1/U1/Z ), .a(\I1/acb ) );
    ao222_1 \I1/U5/U18/U1/U1  ( .x(\I1/ba ), .a(\I1/latch ), .b(n14), .c(
        \I1/latch ), .d(\I1/ba ), .e(n14), .f(\I1/ba ) );
    aoi222_1 \I1/U1664/U28/U30/U1  ( .x(\I1/U1664/x[3] ), .a(\I1/ncd[7] ), .b(
        \I1/ncd[6] ), .c(\I1/ncd[7] ), .d(\I1/U1664/U28/Z ), .e(\I1/ncd[6] ), 
        .f(\I1/U1664/U28/Z ) );
    inv_1 \I1/U1664/U28/U30/Uinv  ( .x(\I1/U1664/U28/Z ), .a(\I1/U1664/x[3] )
         );
    aoi222_1 \I1/U1664/U32/U30/U1  ( .x(\I1/U1664/x[0] ), .a(\I1/ncd[1] ), .b(
        \I1/ncd[0] ), .c(\I1/ncd[1] ), .d(\I1/U1664/U32/Z ), .e(\I1/ncd[0] ), 
        .f(\I1/U1664/U32/Z ) );
    inv_1 \I1/U1664/U32/U30/Uinv  ( .x(\I1/U1664/U32/Z ), .a(\I1/U1664/x[0] )
         );
    aoi222_1 \I1/U1664/U29/U30/U1  ( .x(\I1/U1664/x[2] ), .a(\I1/ncd[5] ), .b(
        \I1/ncd[4] ), .c(\I1/ncd[5] ), .d(\I1/U1664/U29/Z ), .e(\I1/ncd[4] ), 
        .f(\I1/U1664/U29/Z ) );
    inv_1 \I1/U1664/U29/U30/Uinv  ( .x(\I1/U1664/U29/Z ), .a(\I1/U1664/x[2] )
         );
    aoi222_1 \I1/U1664/U33/U30/U1  ( .x(\I1/U1664/y[0] ), .a(\I1/U1664/x[1] ), 
        .b(\I1/U1664/x[0] ), .c(\I1/U1664/x[1] ), .d(\I1/U1664/U33/Z ), .e(
        \I1/U1664/x[0] ), .f(\I1/U1664/U33/Z ) );
    inv_1 \I1/U1664/U33/U30/Uinv  ( .x(\I1/U1664/U33/Z ), .a(\I1/U1664/y[0] )
         );
    aoi222_1 \I1/U1664/U30/U30/U1  ( .x(\I1/U1664/y[1] ), .a(\I1/U1664/x[3] ), 
        .b(\I1/U1664/x[2] ), .c(\I1/U1664/x[3] ), .d(\I1/U1664/U30/Z ), .e(
        \I1/U1664/x[2] ), .f(\I1/U1664/U30/Z ) );
    inv_1 \I1/U1664/U30/U30/Uinv  ( .x(\I1/U1664/U30/Z ), .a(\I1/U1664/y[1] )
         );
    aoi222_1 \I1/U1664/U31/U30/U1  ( .x(\I1/U1664/x[1] ), .a(\I1/ncd[3] ), .b(
        \I1/ncd[2] ), .c(\I1/ncd[3] ), .d(\I1/U1664/U31/Z ), .e(\I1/ncd[2] ), 
        .f(\I1/U1664/U31/Z ) );
    inv_1 \I1/U1664/U31/U30/Uinv  ( .x(\I1/U1664/U31/Z ), .a(\I1/U1664/x[1] )
         );
    aoi222_1 \I1/U1664/U37/U30/U1  ( .x(\I1/localcd ), .a(\I1/U1664/y[0] ), 
        .b(\I1/U1664/y[1] ), .c(\I1/U1664/y[0] ), .d(\I1/U1664/U37/Z ), .e(
        \I1/U1664/y[1] ), .f(\I1/U1664/U37/Z ) );
    inv_1 \I1/U1664/U37/U30/Uinv  ( .x(\I1/U1664/U37/Z ), .a(\I1/localcd ) );
    nor3_1 \I1/U1669/Unr  ( .x(\I1/U1669/nr ), .a(\I1/ctrlack_internal ), .b(
        n4), .c(\I1/drivel ) );
    nand3_1 \I1/U1669/Und  ( .x(\I1/U1669/nd ), .a(\I1/ctrlack_internal ), .b(
        \I1/driveh ), .c(\I1/drivel ) );
    oa21_1 \I1/U1669/U1  ( .x(\I1/U1669/n2 ), .a(\I1/U1669/n2 ), .b(
        \I1/U1669/nr ), .c(\I1/U1669/nd ) );
    inv_2 \I1/U1669/U3  ( .x(read_lhw), .a(\I1/U1669/n2 ) );
    buf_2 \I2/U1653  ( .x(\I2/latch ), .a(net170) );
    nor2_1 \I2/U264/U5  ( .x(\I2/nlocalcd ), .a(reset), .b(\I2/localcd ) );
    nor2_1 \I2/U1659_0_/U5  ( .x(\I2/ncd[0] ), .a(rd[16]), .b(rd[48]) );
    nor2_1 \I2/U1659_1_/U5  ( .x(\I2/ncd[1] ), .a(rd[17]), .b(rd[49]) );
    nor2_1 \I2/U1659_2_/U5  ( .x(\I2/ncd[2] ), .a(rd[18]), .b(rd[50]) );
    nor2_1 \I2/U1659_3_/U5  ( .x(\I2/ncd[3] ), .a(rd[19]), .b(rd[51]) );
    nor2_1 \I2/U1659_4_/U5  ( .x(\I2/ncd[4] ), .a(rd[20]), .b(rd[52]) );
    nor2_1 \I2/U1659_5_/U5  ( .x(\I2/ncd[5] ), .a(rd[21]), .b(rd[53]) );
    nor2_1 \I2/U1659_6_/U5  ( .x(\I2/ncd[6] ), .a(rd[22]), .b(rd[54]) );
    nor2_1 \I2/U1659_7_/U5  ( .x(\I2/ncd[7] ), .a(rd[23]), .b(rd[55]) );
    nor2_1 \I2/U3/U5  ( .x(\I2/ctrlack_internal ), .a(\I2/acb ), .b(\I2/ba )
         );
    buf_2 \I2/U1665/U7  ( .x(\I2/driveh ), .a(net94) );
    buf_2 \I2/U1666/U7  ( .x(\I2/drivel ), .a(net94) );
    ao23_1 \I2/U1658_0_/U21/U1/U1  ( .x(rd[16]), .a(n2), .b(rd[16]), .c(
        \I2/drivel ), .d(cbl[0]), .e(n1) );
    ao23_1 \I2/U1658_1_/U21/U1/U1  ( .x(rd[17]), .a(n2), .b(rd[17]), .c(
        \I2/driveh ), .d(cbl[1]), .e(n1) );
    ao23_1 \I2/U1658_2_/U21/U1/U1  ( .x(rd[18]), .a(\I2/driveh ), .b(rd[18]), 
        .c(n2), .d(cbl[2]), .e(n1) );
    ao23_1 \I2/U1658_3_/U21/U1/U1  ( .x(rd[19]), .a(n2), .b(rd[19]), .c(
        \I2/driveh ), .d(cbl[3]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_4_/U21/U1/U1  ( .x(rd[20]), .a(\I2/drivel ), .b(rd[20]), 
        .c(n2), .d(cbl[4]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_5_/U21/U1/U1  ( .x(rd[21]), .a(\I2/drivel ), .b(rd[21]), 
        .c(n2), .d(cbl[5]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_6_/U21/U1/U1  ( .x(rd[22]), .a(\I2/driveh ), .b(rd[22]), 
        .c(\I2/drivel ), .d(cbl[6]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_7_/U21/U1/U1  ( .x(rd[23]), .a(\I2/driveh ), .b(rd[23]), 
        .c(\I2/driveh ), .d(cbl[7]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_0_/U21/U1/U1  ( .x(rd[48]), .a(\I2/drivel ), .b(rd[48]), 
        .c(n2), .d(cbh[0]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_1_/U21/U1/U1  ( .x(rd[49]), .a(\I2/driveh ), .b(rd[49]), 
        .c(\I2/drivel ), .d(cbh[1]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_2_/U21/U1/U1  ( .x(rd[50]), .a(\I2/drivel ), .b(rd[50]), 
        .c(\I2/drivel ), .d(cbh[2]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_3_/U21/U1/U1  ( .x(rd[51]), .a(\I2/driveh ), .b(rd[51]), 
        .c(\I2/driveh ), .d(cbh[3]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_4_/U21/U1/U1  ( .x(rd[52]), .a(\I2/drivel ), .b(rd[52]), 
        .c(\I2/driveh ), .d(cbh[4]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_5_/U21/U1/U1  ( .x(rd[53]), .a(\I2/driveh ), .b(rd[53]), 
        .c(n2), .d(cbh[5]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_6_/U21/U1/U1  ( .x(rd[54]), .a(n2), .b(rd[54]), .c(
        \I2/drivel ), .d(cbh[6]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_7_/U21/U1/U1  ( .x(rd[55]), .a(n2), .b(rd[55]), .c(n2), 
        .d(cbh[7]), .e(\I2/latch ) );
    aoai211_1 \I2/U4/U28/U1/U1  ( .x(\I2/U4/U28/U1/clr ), .a(net94), .b(
        \I2/acb ), .c(\I2/nlocalcd ), .d(net170) );
    nand3_1 \I2/U4/U28/U1/U2  ( .x(\I2/U4/U28/U1/set ), .a(\I2/nlocalcd ), .b(
        net94), .c(\I2/acb ) );
    nand2_2 \I2/U4/U28/U1/U3  ( .x(net170), .a(\I2/U4/U28/U1/clr ), .b(
        \I2/U4/U28/U1/set ) );
    oai21_1 \I2/U1/U30/U1/U1  ( .x(\I2/acb ), .a(\I2/U1/Z ), .b(\I2/ba ), .c(
        net94) );
    inv_1 \I2/U1/U30/U1/U2  ( .x(\I2/U1/Z ), .a(\I2/acb ) );
    ao222_1 \I2/U5/U18/U1/U1  ( .x(\I2/ba ), .a(\I2/latch ), .b(n14), .c(
        \I2/latch ), .d(\I2/ba ), .e(n14), .f(\I2/ba ) );
    aoi222_1 \I2/U1664/U28/U30/U1  ( .x(\I2/U1664/x[3] ), .a(\I2/ncd[7] ), .b(
        \I2/ncd[6] ), .c(\I2/ncd[7] ), .d(\I2/U1664/U28/Z ), .e(\I2/ncd[6] ), 
        .f(\I2/U1664/U28/Z ) );
    inv_1 \I2/U1664/U28/U30/Uinv  ( .x(\I2/U1664/U28/Z ), .a(\I2/U1664/x[3] )
         );
    aoi222_1 \I2/U1664/U32/U30/U1  ( .x(\I2/U1664/x[0] ), .a(\I2/ncd[1] ), .b(
        \I2/ncd[0] ), .c(\I2/ncd[1] ), .d(\I2/U1664/U32/Z ), .e(\I2/ncd[0] ), 
        .f(\I2/U1664/U32/Z ) );
    inv_1 \I2/U1664/U32/U30/Uinv  ( .x(\I2/U1664/U32/Z ), .a(\I2/U1664/x[0] )
         );
    aoi222_1 \I2/U1664/U29/U30/U1  ( .x(\I2/U1664/x[2] ), .a(\I2/ncd[5] ), .b(
        \I2/ncd[4] ), .c(\I2/ncd[5] ), .d(\I2/U1664/U29/Z ), .e(\I2/ncd[4] ), 
        .f(\I2/U1664/U29/Z ) );
    inv_1 \I2/U1664/U29/U30/Uinv  ( .x(\I2/U1664/U29/Z ), .a(\I2/U1664/x[2] )
         );
    aoi222_1 \I2/U1664/U33/U30/U1  ( .x(\I2/U1664/y[0] ), .a(\I2/U1664/x[1] ), 
        .b(\I2/U1664/x[0] ), .c(\I2/U1664/x[1] ), .d(\I2/U1664/U33/Z ), .e(
        \I2/U1664/x[0] ), .f(\I2/U1664/U33/Z ) );
    inv_1 \I2/U1664/U33/U30/Uinv  ( .x(\I2/U1664/U33/Z ), .a(\I2/U1664/y[0] )
         );
    aoi222_1 \I2/U1664/U30/U30/U1  ( .x(\I2/U1664/y[1] ), .a(\I2/U1664/x[3] ), 
        .b(\I2/U1664/x[2] ), .c(\I2/U1664/x[3] ), .d(\I2/U1664/U30/Z ), .e(
        \I2/U1664/x[2] ), .f(\I2/U1664/U30/Z ) );
    inv_1 \I2/U1664/U30/U30/Uinv  ( .x(\I2/U1664/U30/Z ), .a(\I2/U1664/y[1] )
         );
    aoi222_1 \I2/U1664/U31/U30/U1  ( .x(\I2/U1664/x[1] ), .a(\I2/ncd[3] ), .b(
        \I2/ncd[2] ), .c(\I2/ncd[3] ), .d(\I2/U1664/U31/Z ), .e(\I2/ncd[2] ), 
        .f(\I2/U1664/U31/Z ) );
    inv_1 \I2/U1664/U31/U30/Uinv  ( .x(\I2/U1664/U31/Z ), .a(\I2/U1664/x[1] )
         );
    aoi222_1 \I2/U1664/U37/U30/U1  ( .x(\I2/localcd ), .a(\I2/U1664/y[0] ), 
        .b(\I2/U1664/y[1] ), .c(\I2/U1664/y[0] ), .d(\I2/U1664/U37/Z ), .e(
        \I2/U1664/y[1] ), .f(\I2/U1664/U37/Z ) );
    inv_1 \I2/U1664/U37/U30/Uinv  ( .x(\I2/U1664/U37/Z ), .a(\I2/localcd ) );
    nor3_1 \I2/U1669/Unr  ( .x(\I2/U1669/nr ), .a(\I2/ctrlack_internal ), .b(
        n2), .c(\I2/drivel ) );
    nand3_1 \I2/U1669/Und  ( .x(\I2/U1669/nd ), .a(\I2/ctrlack_internal ), .b(
        \I2/driveh ), .c(\I2/drivel ) );
    oa21_1 \I2/U1669/U1  ( .x(\I2/U1669/n2 ), .a(\I2/U1669/n2 ), .b(
        \I2/U1669/nr ), .c(\I2/U1669/nd ) );
    inv_2 \I2/U1669/U3  ( .x(net103), .a(\I2/U1669/n2 ) );
    buf_1 U1 ( .x(n1), .a(\I2/latch ) );
    buf_2 U2 ( .x(n2), .a(net94) );
    buf_1 U3 ( .x(n3), .a(\I1/latch ) );
    buf_2 U4 ( .x(n4), .a(net103) );
    buf_1 U5 ( .x(n5), .a(\U1666/latch ) );
    buf_2 U6 ( .x(n6), .a(read) );
    buf_1 U7 ( .x(n7), .a(\U1650/latch ) );
    buf_1 U8 ( .x(n8), .a(\U1650/driveh ) );
    buf_1 U9 ( .x(n9), .a(\U1650/drivel ) );
    buf_1 U10 ( .x(n10), .a(\U1667/latch ) );
    buf_2 U11 ( .x(n11), .a(read_lhw) );
    buf_1 U12 ( .x(n12), .a(\I6/latch ) );
    buf_2 U13 ( .x(n13), .a(net139) );
    buf_3 U14 ( .x(n14), .a(bpullcd) );
    buf_3 U15 ( .x(err[0]), .a(n18) );
    buf_3 U16 ( .x(err[1]), .a(n17) );
endmodule


module chain_fr2dr_byte_5 ( nia, oh, ol, i, nReset, noa );
output [7:0] oh;
output [7:0] ol;
input  [4:0] i;
input  nReset, noa;
output nia;
    wire eop, net135, nca, nbReset, ncla, \c[3] , \c[2] , \c[1] , \c[0] , 
        \cl[3] , \cl[2] , \cl[1] , \cl[0] , asel, bsel, asela, bsela, csel, 
        dsel, csela, dsela, esel, fsel, esela, fsela, naa, nda, \a[3] , \a[2] , 
        \a[1] , \a[0] , \d[3] , \d[2] , \d[1] , \d[0] , nba, nea, nfa, \b[3] , 
        \b[2] , \b[1] , \b[0] , \f[3] , \f[2] , \f[1] , \f[0] , \e[3] , \e[2] , 
        \e[1] , \e[0] , \U891/nack , \U891/acka , \U891/naack[0] , 
        \U891/naack[1] , \U891/iay , \U891/ackb , \U891/reset , \U891/neopack , 
        \U891/U1128/nb , \U891/U1128/na , \U891/U1118_0_/nr , 
        \U891/U1118_0_/nd , \U891/U1118_0_/n2 , \U891/U1118_1_/nr , 
        \U891/U1118_1_/nd , \U891/U1118_1_/n2 , \U891/U1118_2_/nr , 
        \U891/U1118_2_/nd , \U891/U1118_2_/n2 , \U891/U1118_3_/nr , 
        \U891/U1118_3_/nd , \U891/U1118_3_/n2 , \U891/U1117_0_/nr , 
        \U891/U1117_0_/nd , \U891/U1117_0_/n2 , \U891/U1117_1_/nr , 
        \U891/U1117_1_/nd , \U891/U1117_1_/n2 , \U891/U1117_2_/nr , 
        \U891/U1117_2_/nd , \U891/U1117_2_/n2 , \U891/U1117_3_/nr , 
        \U891/U1117_3_/nd , \U891/U1117_3_/n2 , \U886/nack , \U886/acka , 
        \U886/ackb , \U886/reset , \U886/U1128/nb , \U886/U1128/na , 
        \U886/U1127/n5 , \U886/U1127/n1 , \U886/U1127/n2 , \U886/U1127/n3 , 
        \U886/U1127/n4 , \U886/U1118_0_/nr , \U886/U1118_0_/nd , 
        \U886/U1118_0_/n2 , \U886/U1118_1_/nr , \U886/U1118_1_/nd , 
        \U886/U1118_1_/n2 , \U886/U1118_2_/nr , \U886/U1118_2_/nd , 
        \U886/U1118_2_/n2 , \U886/U1118_3_/nr , \U886/U1118_3_/nd , 
        \U886/U1118_3_/n2 , \U886/U1117_0_/nr , \U886/U1117_0_/nd , 
        \U886/U1117_0_/n2 , \U886/U1117_1_/nr , \U886/U1117_1_/nd , 
        \U886/U1117_1_/n2 , \U886/U1117_2_/nr , \U886/U1117_2_/nd , 
        \U886/U1117_2_/n2 , \U886/U1117_3_/nr , \U886/U1117_3_/nd , 
        \U886/U1117_3_/n2 , \U884/nack , \U884/acka , \U884/ackb , 
        \U884/reset , \U884/U1128/nb , \U884/U1128/na , \U884/U1127/n5 , 
        \U884/U1127/n1 , \U884/U1127/n2 , \U884/U1127/n3 , \U884/U1127/n4 , 
        \U884/U1118_0_/nr , \U884/U1118_0_/nd , \U884/U1118_0_/n2 , 
        \U884/U1118_1_/nr , \U884/U1118_1_/nd , \U884/U1118_1_/n2 , 
        \U884/U1118_2_/nr , \U884/U1118_2_/nd , \U884/U1118_2_/n2 , 
        \U884/U1118_3_/nr , \U884/U1118_3_/nd , \U884/U1118_3_/n2 , 
        \U884/U1117_0_/nr , \U884/U1117_0_/nd , \U884/U1117_0_/n2 , 
        \U884/U1117_1_/nr , \U884/U1117_1_/nd , \U884/U1117_1_/n2 , 
        \U884/U1117_2_/nr , \U884/U1117_2_/nd , \U884/U1117_2_/n2 , 
        \U884/U1117_3_/nr , \U884/U1117_3_/nd , \U884/U1117_3_/n2 , 
        \U888/naack , \U888/r , \U888/s , \U888/nback , \U888/reset , 
        \U887/naack , \U887/r , \U887/s , \U887/nback , \U887/reset , 
        \U885/naack , \U885/r , \U885/s , \U885/nback , \U885/reset , \U877/x , 
        \U877/y , \U877/reset , \U877/U590/U25/U1/clr , \U877/U590/U25/U1/ob , 
        \U877/U589/U25/U1/clr , \U877/U589/U25/U1/ob , \U877/U588/U25/U1/clr , 
        \U877/U588/U25/U1/ob , \U877/U591/U25/U1/clr , \U877/U591/U25/U1/ob , 
        \U876/x , \U876/y , \U876/reset , \U876/U590/U25/U1/clr , 
        \U876/U590/U25/U1/ob , \U876/U589/U25/U1/clr , \U876/U589/U25/U1/ob , 
        \U876/U588/U25/U1/clr , \U876/U588/U25/U1/ob , \U876/U591/U25/U1/clr , 
        \U876/U591/U25/U1/ob , \U2/x , \U2/y , \U2/reset , 
        \U2/U590/U25/U1/clr , \U2/U590/U25/U1/ob , \U2/U589/U25/U1/clr , 
        \U2/U589/U25/U1/ob , \U2/U588/U25/U1/clr , \U2/U588/U25/U1/ob , 
        \U2/U591/U25/U1/clr , \U2/U591/U25/U1/ob , \U1/x , \U1/y , \U1/reset , 
        \U1/U590/U25/U1/clr , \U1/U590/U25/U1/ob , \U1/U589/U25/U1/clr , 
        \U1/U589/U25/U1/ob , \U1/U588/U25/U1/clr , \U1/U588/U25/U1/ob , 
        \U1/U591/U25/U1/clr , \U1/U591/U25/U1/ob , \U881/nack[1] , 
        \U881/nack[0] , n1;
    buf_2 U897 ( .x(nbReset), .a(nReset) );
    and4_1 \U894/U12  ( .x(eop), .a(ncla), .b(csela), .c(asela), .d(i[4]) );
    inv_1 \U891/U1126/U3  ( .x(\U891/reset ), .a(nbReset) );
    inv_1 \U891/U1139/U3  ( .x(\U891/neopack ), .a(eop) );
    nand3_1 \U891/U1131/U9  ( .x(\U891/iay ), .a(\U891/neopack ), .b(
        \U891/naack[0] ), .c(\U891/naack[1] ) );
    nor3_1 \U891/U1128/U27  ( .x(\U891/U1128/nb ), .a(\U891/reset ), .b(\b[3] 
        ), .c(\b[2] ) );
    nor2_1 \U891/U1128/U26  ( .x(\U891/U1128/na ), .a(\b[1] ), .b(\b[0] ) );
    nand2_2 \U891/U1128/U29  ( .x(\U891/ackb ), .a(\U891/U1128/nb ), .b(
        \U891/U1128/na ) );
    nor2_1 \U891/U1133/U5  ( .x(\U891/naack[0] ), .a(\a[3] ), .b(\a[2] ) );
    nor2_1 \U891/U1108/U5  ( .x(\U891/nack ), .a(\U891/acka ), .b(\U891/ackb )
         );
    nor2_1 \U891/U1134/U5  ( .x(\U891/naack[1] ), .a(\a[1] ), .b(\a[0] ) );
    nor2_2 \U891/U914/U6  ( .x(nia), .a(\U891/iay ), .b(\U891/ackb ) );
    nand2_1 \U891/U1130/U5  ( .x(\U891/acka ), .a(\U891/naack[0] ), .b(
        \U891/naack[1] ) );
    ao222_4 \U891/U1121/U1/U1  ( .x(bsela), .a(\U891/nack ), .b(bsel), .c(
        \U891/nack ), .d(bsela), .e(bsel), .f(bsela) );
    ao222_4 \U891/U1120/U1/U1  ( .x(asela), .a(asel), .b(\U891/nack ), .c(asel
        ), .d(asela), .e(\U891/nack ), .f(asela) );
    nor3_1 \U891/U1118_0_/Unr  ( .x(\U891/U1118_0_/nr ), .a(i[0]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_0_/Und  ( .x(\U891/U1118_0_/nd ), .a(i[0]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_0_/U1  ( .x(\U891/U1118_0_/n2 ), .a(\U891/U1118_0_/n2 ), 
        .b(\U891/U1118_0_/nr ), .c(\U891/U1118_0_/nd ) );
    inv_2 \U891/U1118_0_/U3  ( .x(\a[0] ), .a(\U891/U1118_0_/n2 ) );
    nor3_1 \U891/U1118_1_/Unr  ( .x(\U891/U1118_1_/nr ), .a(i[1]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_1_/Und  ( .x(\U891/U1118_1_/nd ), .a(i[1]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_1_/U1  ( .x(\U891/U1118_1_/n2 ), .a(\U891/U1118_1_/n2 ), 
        .b(\U891/U1118_1_/nr ), .c(\U891/U1118_1_/nd ) );
    inv_2 \U891/U1118_1_/U3  ( .x(\a[1] ), .a(\U891/U1118_1_/n2 ) );
    nor3_1 \U891/U1118_2_/Unr  ( .x(\U891/U1118_2_/nr ), .a(i[2]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_2_/Und  ( .x(\U891/U1118_2_/nd ), .a(i[2]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_2_/U1  ( .x(\U891/U1118_2_/n2 ), .a(\U891/U1118_2_/n2 ), 
        .b(\U891/U1118_2_/nr ), .c(\U891/U1118_2_/nd ) );
    inv_2 \U891/U1118_2_/U3  ( .x(\a[2] ), .a(\U891/U1118_2_/n2 ) );
    nor3_1 \U891/U1118_3_/Unr  ( .x(\U891/U1118_3_/nr ), .a(i[3]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_3_/Und  ( .x(\U891/U1118_3_/nd ), .a(i[3]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_3_/U1  ( .x(\U891/U1118_3_/n2 ), .a(\U891/U1118_3_/n2 ), 
        .b(\U891/U1118_3_/nr ), .c(\U891/U1118_3_/nd ) );
    inv_2 \U891/U1118_3_/U3  ( .x(\a[3] ), .a(\U891/U1118_3_/n2 ) );
    nor3_1 \U891/U1117_0_/Unr  ( .x(\U891/U1117_0_/nr ), .a(i[0]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_0_/Und  ( .x(\U891/U1117_0_/nd ), .a(i[0]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_0_/U1  ( .x(\U891/U1117_0_/n2 ), .a(\U891/U1117_0_/n2 ), 
        .b(\U891/U1117_0_/nr ), .c(\U891/U1117_0_/nd ) );
    inv_2 \U891/U1117_0_/U3  ( .x(\b[0] ), .a(\U891/U1117_0_/n2 ) );
    nor3_1 \U891/U1117_1_/Unr  ( .x(\U891/U1117_1_/nr ), .a(i[1]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_1_/Und  ( .x(\U891/U1117_1_/nd ), .a(i[1]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_1_/U1  ( .x(\U891/U1117_1_/n2 ), .a(\U891/U1117_1_/n2 ), 
        .b(\U891/U1117_1_/nr ), .c(\U891/U1117_1_/nd ) );
    inv_2 \U891/U1117_1_/U3  ( .x(\b[1] ), .a(\U891/U1117_1_/n2 ) );
    nor3_1 \U891/U1117_2_/Unr  ( .x(\U891/U1117_2_/nr ), .a(i[2]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_2_/Und  ( .x(\U891/U1117_2_/nd ), .a(i[2]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_2_/U1  ( .x(\U891/U1117_2_/n2 ), .a(\U891/U1117_2_/n2 ), 
        .b(\U891/U1117_2_/nr ), .c(\U891/U1117_2_/nd ) );
    inv_2 \U891/U1117_2_/U3  ( .x(\b[2] ), .a(\U891/U1117_2_/n2 ) );
    nor3_1 \U891/U1117_3_/Unr  ( .x(\U891/U1117_3_/nr ), .a(i[3]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_3_/Und  ( .x(\U891/U1117_3_/nd ), .a(i[3]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_3_/U1  ( .x(\U891/U1117_3_/n2 ), .a(\U891/U1117_3_/n2 ), 
        .b(\U891/U1117_3_/nr ), .c(\U891/U1117_3_/nd ) );
    inv_2 \U891/U1117_3_/U3  ( .x(\b[3] ), .a(\U891/U1117_3_/n2 ) );
    inv_1 \U886/U1126/U3  ( .x(\U886/reset ), .a(nbReset) );
    nor3_1 \U886/U1128/U27  ( .x(\U886/U1128/nb ), .a(\U886/reset ), .b(\f[3] 
        ), .c(\f[2] ) );
    nor2_1 \U886/U1128/U26  ( .x(\U886/U1128/na ), .a(\f[1] ), .b(\f[0] ) );
    nand2_2 \U886/U1128/U29  ( .x(\U886/ackb ), .a(\U886/U1128/nb ), .b(
        \U886/U1128/na ) );
    nor2_1 \U886/U1108/U5  ( .x(\U886/nack ), .a(\U886/acka ), .b(\U886/ackb )
         );
    nor2_2 \U886/U914/U6  ( .x(nba), .a(\U886/acka ), .b(\U886/ackb ) );
    and4_1 \U886/U1127/U25  ( .x(\U886/U1127/n5 ), .a(\U886/U1127/n1 ), .b(
        \U886/U1127/n2 ), .c(\U886/U1127/n3 ), .d(\U886/U1127/n4 ) );
    inv_1 \U886/U1127/U1  ( .x(\U886/U1127/n1 ), .a(\e[3] ) );
    inv_1 \U886/U1127/U2  ( .x(\U886/U1127/n2 ), .a(\e[2] ) );
    inv_1 \U886/U1127/U3  ( .x(\U886/U1127/n3 ), .a(\e[1] ) );
    inv_1 \U886/U1127/U4  ( .x(\U886/U1127/n4 ), .a(\e[0] ) );
    inv_2 \U886/U1127/U5  ( .x(\U886/acka ), .a(\U886/U1127/n5 ) );
    ao222_2 \U886/U1121/U19/U1/U1  ( .x(fsela), .a(\U886/nack ), .b(fsel), .c(
        \U886/nack ), .d(fsela), .e(fsel), .f(fsela) );
    ao222_2 \U886/U1120/U19/U1/U1  ( .x(esela), .a(esel), .b(\U886/nack ), .c(
        esel), .d(esela), .e(\U886/nack ), .f(esela) );
    nor3_1 \U886/U1118_0_/Unr  ( .x(\U886/U1118_0_/nr ), .a(\b[0] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_0_/Und  ( .x(\U886/U1118_0_/nd ), .a(\b[0] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_0_/U1  ( .x(\U886/U1118_0_/n2 ), .a(\U886/U1118_0_/n2 ), 
        .b(\U886/U1118_0_/nr ), .c(\U886/U1118_0_/nd ) );
    inv_2 \U886/U1118_0_/U3  ( .x(\e[0] ), .a(\U886/U1118_0_/n2 ) );
    nor3_1 \U886/U1118_1_/Unr  ( .x(\U886/U1118_1_/nr ), .a(\b[1] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_1_/Und  ( .x(\U886/U1118_1_/nd ), .a(\b[1] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_1_/U1  ( .x(\U886/U1118_1_/n2 ), .a(\U886/U1118_1_/n2 ), 
        .b(\U886/U1118_1_/nr ), .c(\U886/U1118_1_/nd ) );
    inv_2 \U886/U1118_1_/U3  ( .x(\e[1] ), .a(\U886/U1118_1_/n2 ) );
    nor3_1 \U886/U1118_2_/Unr  ( .x(\U886/U1118_2_/nr ), .a(\b[2] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_2_/Und  ( .x(\U886/U1118_2_/nd ), .a(\b[2] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_2_/U1  ( .x(\U886/U1118_2_/n2 ), .a(\U886/U1118_2_/n2 ), 
        .b(\U886/U1118_2_/nr ), .c(\U886/U1118_2_/nd ) );
    inv_2 \U886/U1118_2_/U3  ( .x(\e[2] ), .a(\U886/U1118_2_/n2 ) );
    nor3_1 \U886/U1118_3_/Unr  ( .x(\U886/U1118_3_/nr ), .a(\b[3] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_3_/Und  ( .x(\U886/U1118_3_/nd ), .a(\b[3] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_3_/U1  ( .x(\U886/U1118_3_/n2 ), .a(\U886/U1118_3_/n2 ), 
        .b(\U886/U1118_3_/nr ), .c(\U886/U1118_3_/nd ) );
    inv_2 \U886/U1118_3_/U3  ( .x(\e[3] ), .a(\U886/U1118_3_/n2 ) );
    nor3_1 \U886/U1117_0_/Unr  ( .x(\U886/U1117_0_/nr ), .a(\b[0] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_0_/Und  ( .x(\U886/U1117_0_/nd ), .a(\b[0] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_0_/U1  ( .x(\U886/U1117_0_/n2 ), .a(\U886/U1117_0_/n2 ), 
        .b(\U886/U1117_0_/nr ), .c(\U886/U1117_0_/nd ) );
    inv_2 \U886/U1117_0_/U3  ( .x(\f[0] ), .a(\U886/U1117_0_/n2 ) );
    nor3_1 \U886/U1117_1_/Unr  ( .x(\U886/U1117_1_/nr ), .a(\b[1] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_1_/Und  ( .x(\U886/U1117_1_/nd ), .a(\b[1] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_1_/U1  ( .x(\U886/U1117_1_/n2 ), .a(\U886/U1117_1_/n2 ), 
        .b(\U886/U1117_1_/nr ), .c(\U886/U1117_1_/nd ) );
    inv_2 \U886/U1117_1_/U3  ( .x(\f[1] ), .a(\U886/U1117_1_/n2 ) );
    nor3_1 \U886/U1117_2_/Unr  ( .x(\U886/U1117_2_/nr ), .a(\b[2] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_2_/Und  ( .x(\U886/U1117_2_/nd ), .a(\b[2] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_2_/U1  ( .x(\U886/U1117_2_/n2 ), .a(\U886/U1117_2_/n2 ), 
        .b(\U886/U1117_2_/nr ), .c(\U886/U1117_2_/nd ) );
    inv_2 \U886/U1117_2_/U3  ( .x(\f[2] ), .a(\U886/U1117_2_/n2 ) );
    nor3_1 \U886/U1117_3_/Unr  ( .x(\U886/U1117_3_/nr ), .a(\b[3] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_3_/Und  ( .x(\U886/U1117_3_/nd ), .a(\b[3] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_3_/U1  ( .x(\U886/U1117_3_/n2 ), .a(\U886/U1117_3_/n2 ), 
        .b(\U886/U1117_3_/nr ), .c(\U886/U1117_3_/nd ) );
    inv_2 \U886/U1117_3_/U3  ( .x(\f[3] ), .a(\U886/U1117_3_/n2 ) );
    inv_1 \U884/U1126/U3  ( .x(\U884/reset ), .a(nbReset) );
    nor3_1 \U884/U1128/U27  ( .x(\U884/U1128/nb ), .a(\U884/reset ), .b(\d[3] 
        ), .c(\d[2] ) );
    nor2_1 \U884/U1128/U26  ( .x(\U884/U1128/na ), .a(\d[1] ), .b(\d[0] ) );
    nand2_2 \U884/U1128/U29  ( .x(\U884/ackb ), .a(\U884/U1128/nb ), .b(
        \U884/U1128/na ) );
    nor2_1 \U884/U1108/U5  ( .x(\U884/nack ), .a(\U884/acka ), .b(\U884/ackb )
         );
    nor2_2 \U884/U914/U6  ( .x(naa), .a(\U884/acka ), .b(\U884/ackb ) );
    and4_1 \U884/U1127/U25  ( .x(\U884/U1127/n5 ), .a(\U884/U1127/n1 ), .b(
        \U884/U1127/n2 ), .c(\U884/U1127/n3 ), .d(\U884/U1127/n4 ) );
    inv_1 \U884/U1127/U1  ( .x(\U884/U1127/n1 ), .a(\c[3] ) );
    inv_1 \U884/U1127/U2  ( .x(\U884/U1127/n2 ), .a(\c[2] ) );
    inv_1 \U884/U1127/U3  ( .x(\U884/U1127/n3 ), .a(\c[1] ) );
    inv_1 \U884/U1127/U4  ( .x(\U884/U1127/n4 ), .a(\c[0] ) );
    inv_2 \U884/U1127/U5  ( .x(\U884/acka ), .a(\U884/U1127/n5 ) );
    ao222_2 \U884/U1121/U19/U1/U1  ( .x(dsela), .a(\U884/nack ), .b(dsel), .c(
        \U884/nack ), .d(dsela), .e(dsel), .f(dsela) );
    ao222_2 \U884/U1120/U19/U1/U1  ( .x(csela), .a(csel), .b(\U884/nack ), .c(
        csel), .d(csela), .e(\U884/nack ), .f(csela) );
    nor3_1 \U884/U1118_0_/Unr  ( .x(\U884/U1118_0_/nr ), .a(\a[0] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_0_/Und  ( .x(\U884/U1118_0_/nd ), .a(\a[0] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_0_/U1  ( .x(\U884/U1118_0_/n2 ), .a(\U884/U1118_0_/n2 ), 
        .b(\U884/U1118_0_/nr ), .c(\U884/U1118_0_/nd ) );
    inv_2 \U884/U1118_0_/U3  ( .x(\c[0] ), .a(\U884/U1118_0_/n2 ) );
    nor3_1 \U884/U1118_1_/Unr  ( .x(\U884/U1118_1_/nr ), .a(\a[1] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_1_/Und  ( .x(\U884/U1118_1_/nd ), .a(\a[1] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_1_/U1  ( .x(\U884/U1118_1_/n2 ), .a(\U884/U1118_1_/n2 ), 
        .b(\U884/U1118_1_/nr ), .c(\U884/U1118_1_/nd ) );
    inv_2 \U884/U1118_1_/U3  ( .x(\c[1] ), .a(\U884/U1118_1_/n2 ) );
    nor3_1 \U884/U1118_2_/Unr  ( .x(\U884/U1118_2_/nr ), .a(\a[2] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_2_/Und  ( .x(\U884/U1118_2_/nd ), .a(\a[2] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_2_/U1  ( .x(\U884/U1118_2_/n2 ), .a(\U884/U1118_2_/n2 ), 
        .b(\U884/U1118_2_/nr ), .c(\U884/U1118_2_/nd ) );
    inv_2 \U884/U1118_2_/U3  ( .x(\c[2] ), .a(\U884/U1118_2_/n2 ) );
    nor3_1 \U884/U1118_3_/Unr  ( .x(\U884/U1118_3_/nr ), .a(\a[3] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_3_/Und  ( .x(\U884/U1118_3_/nd ), .a(\a[3] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_3_/U1  ( .x(\U884/U1118_3_/n2 ), .a(\U884/U1118_3_/n2 ), 
        .b(\U884/U1118_3_/nr ), .c(\U884/U1118_3_/nd ) );
    inv_2 \U884/U1118_3_/U3  ( .x(\c[3] ), .a(\U884/U1118_3_/n2 ) );
    nor3_1 \U884/U1117_0_/Unr  ( .x(\U884/U1117_0_/nr ), .a(\a[0] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_0_/Und  ( .x(\U884/U1117_0_/nd ), .a(\a[0] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_0_/U1  ( .x(\U884/U1117_0_/n2 ), .a(\U884/U1117_0_/n2 ), 
        .b(\U884/U1117_0_/nr ), .c(\U884/U1117_0_/nd ) );
    inv_2 \U884/U1117_0_/U3  ( .x(\d[0] ), .a(\U884/U1117_0_/n2 ) );
    nor3_1 \U884/U1117_1_/Unr  ( .x(\U884/U1117_1_/nr ), .a(\a[1] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_1_/Und  ( .x(\U884/U1117_1_/nd ), .a(\a[1] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_1_/U1  ( .x(\U884/U1117_1_/n2 ), .a(\U884/U1117_1_/n2 ), 
        .b(\U884/U1117_1_/nr ), .c(\U884/U1117_1_/nd ) );
    inv_2 \U884/U1117_1_/U3  ( .x(\d[1] ), .a(\U884/U1117_1_/n2 ) );
    nor3_1 \U884/U1117_2_/Unr  ( .x(\U884/U1117_2_/nr ), .a(\a[2] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_2_/Und  ( .x(\U884/U1117_2_/nd ), .a(\a[2] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_2_/U1  ( .x(\U884/U1117_2_/n2 ), .a(\U884/U1117_2_/n2 ), 
        .b(\U884/U1117_2_/nr ), .c(\U884/U1117_2_/nd ) );
    inv_2 \U884/U1117_2_/U3  ( .x(\d[2] ), .a(\U884/U1117_2_/n2 ) );
    nor3_1 \U884/U1117_3_/Unr  ( .x(\U884/U1117_3_/nr ), .a(\a[3] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_3_/Und  ( .x(\U884/U1117_3_/nd ), .a(\a[3] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_3_/U1  ( .x(\U884/U1117_3_/n2 ), .a(\U884/U1117_3_/n2 ), 
        .b(\U884/U1117_3_/nr ), .c(\U884/U1117_3_/nd ) );
    inv_2 \U884/U1117_3_/U3  ( .x(\d[3] ), .a(\U884/U1117_3_/n2 ) );
    nand2_1 \U888/U1128/U5  ( .x(\U888/s ), .a(\U888/r ), .b(\U888/nback ) );
    nand2_1 \U888/U1103/U5  ( .x(\U888/r ), .a(\U888/naack ), .b(\U888/s ) );
    inv_1 \U888/U1111/U3  ( .x(\U888/reset ), .a(nbReset) );
    inv_1 \U888/U1112/U3  ( .x(\U888/naack ), .a(esela) );
    nor2_1 \U888/U1127/U5  ( .x(\U888/nback ), .a(fsela), .b(\U888/reset ) );
    and2_2 \U888/U1129/U8  ( .x(esel), .a(\U888/nback ), .b(\U888/s ) );
    and2_2 \U888/U1124/U8  ( .x(fsel), .a(\U888/r ), .b(\U888/naack ) );
    nand2_1 \U887/U1128/U5  ( .x(\U887/s ), .a(\U887/r ), .b(\U887/nback ) );
    nand2_1 \U887/U1103/U5  ( .x(\U887/r ), .a(\U887/naack ), .b(\U887/s ) );
    inv_1 \U887/U1111/U3  ( .x(\U887/reset ), .a(nbReset) );
    inv_1 \U887/U1112/U3  ( .x(\U887/naack ), .a(csela) );
    nor2_1 \U887/U1127/U5  ( .x(\U887/nback ), .a(dsela), .b(\U887/reset ) );
    and2_2 \U887/U1129/U8  ( .x(csel), .a(\U887/nback ), .b(\U887/s ) );
    and2_2 \U887/U1124/U8  ( .x(dsel), .a(\U887/r ), .b(\U887/naack ) );
    nand2_1 \U885/U1128/U5  ( .x(\U885/s ), .a(\U885/r ), .b(\U885/nback ) );
    nand2_1 \U885/U1103/U5  ( .x(\U885/r ), .a(\U885/naack ), .b(\U885/s ) );
    inv_1 \U885/U1111/U3  ( .x(\U885/reset ), .a(nbReset) );
    inv_1 \U885/U1112/U3  ( .x(\U885/naack ), .a(asela) );
    nor2_1 \U885/U1127/U5  ( .x(\U885/nback ), .a(bsela), .b(\U885/reset ) );
    and2_2 \U885/U1129/U8  ( .x(asel), .a(\U885/nback ), .b(\U885/s ) );
    and2_2 \U885/U1124/U8  ( .x(bsel), .a(\U885/r ), .b(\U885/naack ) );
    nor3_1 \U877/U594/U7  ( .x(\U877/x ), .a(ol[7]), .b(\U877/reset ), .c(oh
        [7]) );
    nor3_1 \U877/U593/U7  ( .x(\U877/y ), .a(ol[6]), .b(\U877/reset ), .c(oh
        [6]) );
    inv_1 \U877/U604/U3  ( .x(\U877/reset ), .a(nbReset) );
    oa31_1 \U877/U590/U25/U1/Uclr  ( .x(\U877/U590/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[1] ), .d(oh[6]) );
    oaoi211_1 \U877/U590/U25/U1/Uaoi  ( .x(\U877/U590/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[1] ), .c(n1), .d(\U877/U590/U25/U1/clr ) );
    inv_2 \U877/U590/U25/U1/Ui  ( .x(oh[6]), .a(\U877/U590/U25/U1/ob ) );
    oa31_1 \U877/U589/U25/U1/Uclr  ( .x(\U877/U589/U25/U1/clr ), .a(net135), 
        .b(\cl[1] ), .c(\cl[0] ), .d(ol[7]) );
    oaoi211_1 \U877/U589/U25/U1/Uaoi  ( .x(\U877/U589/U25/U1/ob ), .a(\cl[1] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U589/U25/U1/clr ) );
    inv_2 \U877/U589/U25/U1/Ui  ( .x(ol[7]), .a(\U877/U589/U25/U1/ob ) );
    oa31_1 \U877/U588/U25/U1/Uclr  ( .x(\U877/U588/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[2] ), .d(oh[7]) );
    oaoi211_1 \U877/U588/U25/U1/Uaoi  ( .x(\U877/U588/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[2] ), .c(n1), .d(\U877/U588/U25/U1/clr ) );
    inv_2 \U877/U588/U25/U1/Ui  ( .x(oh[7]), .a(\U877/U588/U25/U1/ob ) );
    oa31_1 \U877/U591/U25/U1/Uclr  ( .x(\U877/U591/U25/U1/clr ), .a(net135), 
        .b(\cl[2] ), .c(\cl[0] ), .d(ol[6]) );
    oaoi211_1 \U877/U591/U25/U1/Uaoi  ( .x(\U877/U591/U25/U1/ob ), .a(\cl[2] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U591/U25/U1/clr ) );
    inv_2 \U877/U591/U25/U1/Ui  ( .x(ol[6]), .a(\U877/U591/U25/U1/ob ) );
    ao222_2 \U877/U592/U19/U1/U1  ( .x(ncla), .a(\U877/x ), .b(\U877/y ), .c(
        \U877/x ), .d(ncla), .e(\U877/y ), .f(ncla) );
    nor3_1 \U876/U594/U7  ( .x(\U876/x ), .a(ol[3]), .b(\U876/reset ), .c(oh
        [3]) );
    nor3_1 \U876/U593/U7  ( .x(\U876/y ), .a(ol[2]), .b(\U876/reset ), .c(oh
        [2]) );
    inv_1 \U876/U604/U3  ( .x(\U876/reset ), .a(nbReset) );
    oa31_1 \U876/U590/U25/U1/Uclr  ( .x(\U876/U590/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[1] ), .d(oh[2]) );
    oaoi211_1 \U876/U590/U25/U1/Uaoi  ( .x(\U876/U590/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[1] ), .c(n1), .d(\U876/U590/U25/U1/clr ) );
    inv_2 \U876/U590/U25/U1/Ui  ( .x(oh[2]), .a(\U876/U590/U25/U1/ob ) );
    oa31_1 \U876/U589/U25/U1/Uclr  ( .x(\U876/U589/U25/U1/clr ), .a(net135), 
        .b(\d[1] ), .c(\d[0] ), .d(ol[3]) );
    oaoi211_1 \U876/U589/U25/U1/Uaoi  ( .x(\U876/U589/U25/U1/ob ), .a(\d[1] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U589/U25/U1/clr ) );
    inv_2 \U876/U589/U25/U1/Ui  ( .x(ol[3]), .a(\U876/U589/U25/U1/ob ) );
    oa31_1 \U876/U588/U25/U1/Uclr  ( .x(\U876/U588/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[2] ), .d(oh[3]) );
    oaoi211_1 \U876/U588/U25/U1/Uaoi  ( .x(\U876/U588/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[2] ), .c(n1), .d(\U876/U588/U25/U1/clr ) );
    inv_2 \U876/U588/U25/U1/Ui  ( .x(oh[3]), .a(\U876/U588/U25/U1/ob ) );
    oa31_1 \U876/U591/U25/U1/Uclr  ( .x(\U876/U591/U25/U1/clr ), .a(net135), 
        .b(\d[2] ), .c(\d[0] ), .d(ol[2]) );
    oaoi211_1 \U876/U591/U25/U1/Uaoi  ( .x(\U876/U591/U25/U1/ob ), .a(\d[2] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U591/U25/U1/clr ) );
    inv_2 \U876/U591/U25/U1/Ui  ( .x(ol[2]), .a(\U876/U591/U25/U1/ob ) );
    ao222_2 \U876/U592/U19/U1/U1  ( .x(nda), .a(\U876/x ), .b(\U876/y ), .c(
        \U876/x ), .d(nda), .e(\U876/y ), .f(nda) );
    nor3_1 \U2/U594/U7  ( .x(\U2/x ), .a(ol[1]), .b(\U2/reset ), .c(oh[1]) );
    nor3_1 \U2/U593/U7  ( .x(\U2/y ), .a(ol[0]), .b(\U2/reset ), .c(oh[0]) );
    inv_1 \U2/U604/U3  ( .x(\U2/reset ), .a(nbReset) );
    oa31_1 \U2/U590/U25/U1/Uclr  ( .x(\U2/U590/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[1] ), .d(oh[0]) );
    oaoi211_1 \U2/U590/U25/U1/Uaoi  ( .x(\U2/U590/U25/U1/ob ), .a(\f[3] ), .b(
        \f[1] ), .c(n1), .d(\U2/U590/U25/U1/clr ) );
    inv_2 \U2/U590/U25/U1/Ui  ( .x(oh[0]), .a(\U2/U590/U25/U1/ob ) );
    oa31_1 \U2/U589/U25/U1/Uclr  ( .x(\U2/U589/U25/U1/clr ), .a(net135), .b(
        \f[1] ), .c(\f[0] ), .d(ol[1]) );
    oaoi211_1 \U2/U589/U25/U1/Uaoi  ( .x(\U2/U589/U25/U1/ob ), .a(\f[1] ), .b(
        \f[0] ), .c(n1), .d(\U2/U589/U25/U1/clr ) );
    inv_2 \U2/U589/U25/U1/Ui  ( .x(ol[1]), .a(\U2/U589/U25/U1/ob ) );
    oa31_1 \U2/U588/U25/U1/Uclr  ( .x(\U2/U588/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[2] ), .d(oh[1]) );
    oaoi211_1 \U2/U588/U25/U1/Uaoi  ( .x(\U2/U588/U25/U1/ob ), .a(\f[3] ), .b(
        \f[2] ), .c(n1), .d(\U2/U588/U25/U1/clr ) );
    inv_2 \U2/U588/U25/U1/Ui  ( .x(oh[1]), .a(\U2/U588/U25/U1/ob ) );
    oa31_1 \U2/U591/U25/U1/Uclr  ( .x(\U2/U591/U25/U1/clr ), .a(net135), .b(
        \f[2] ), .c(\f[0] ), .d(ol[0]) );
    oaoi211_1 \U2/U591/U25/U1/Uaoi  ( .x(\U2/U591/U25/U1/ob ), .a(\f[2] ), .b(
        \f[0] ), .c(n1), .d(\U2/U591/U25/U1/clr ) );
    inv_2 \U2/U591/U25/U1/Ui  ( .x(ol[0]), .a(\U2/U591/U25/U1/ob ) );
    ao222_2 \U2/U592/U19/U1/U1  ( .x(nfa), .a(\U2/x ), .b(\U2/y ), .c(\U2/x ), 
        .d(nfa), .e(\U2/y ), .f(nfa) );
    nor3_1 \U1/U594/U7  ( .x(\U1/x ), .a(ol[5]), .b(\U1/reset ), .c(oh[5]) );
    nor3_1 \U1/U593/U7  ( .x(\U1/y ), .a(ol[4]), .b(\U1/reset ), .c(oh[4]) );
    inv_1 \U1/U604/U3  ( .x(\U1/reset ), .a(nbReset) );
    oa31_1 \U1/U590/U25/U1/Uclr  ( .x(\U1/U590/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[1] ), .d(oh[4]) );
    oaoi211_1 \U1/U590/U25/U1/Uaoi  ( .x(\U1/U590/U25/U1/ob ), .a(\e[3] ), .b(
        \e[1] ), .c(n1), .d(\U1/U590/U25/U1/clr ) );
    inv_2 \U1/U590/U25/U1/Ui  ( .x(oh[4]), .a(\U1/U590/U25/U1/ob ) );
    oa31_1 \U1/U589/U25/U1/Uclr  ( .x(\U1/U589/U25/U1/clr ), .a(net135), .b(
        \e[1] ), .c(\e[0] ), .d(ol[5]) );
    oaoi211_1 \U1/U589/U25/U1/Uaoi  ( .x(\U1/U589/U25/U1/ob ), .a(\e[1] ), .b(
        \e[0] ), .c(n1), .d(\U1/U589/U25/U1/clr ) );
    inv_2 \U1/U589/U25/U1/Ui  ( .x(ol[5]), .a(\U1/U589/U25/U1/ob ) );
    oa31_1 \U1/U588/U25/U1/Uclr  ( .x(\U1/U588/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[2] ), .d(oh[5]) );
    oaoi211_1 \U1/U588/U25/U1/Uaoi  ( .x(\U1/U588/U25/U1/ob ), .a(\e[3] ), .b(
        \e[2] ), .c(n1), .d(\U1/U588/U25/U1/clr ) );
    inv_2 \U1/U588/U25/U1/Ui  ( .x(oh[5]), .a(\U1/U588/U25/U1/ob ) );
    oa31_1 \U1/U591/U25/U1/Uclr  ( .x(\U1/U591/U25/U1/clr ), .a(net135), .b(
        \e[2] ), .c(\e[0] ), .d(ol[4]) );
    oaoi211_1 \U1/U591/U25/U1/Uaoi  ( .x(\U1/U591/U25/U1/ob ), .a(\e[2] ), .b(
        \e[0] ), .c(n1), .d(\U1/U591/U25/U1/clr ) );
    inv_2 \U1/U591/U25/U1/Ui  ( .x(ol[4]), .a(\U1/U591/U25/U1/ob ) );
    ao222_2 \U1/U592/U19/U1/U1  ( .x(nea), .a(\U1/x ), .b(\U1/y ), .c(\U1/x ), 
        .d(nea), .e(\U1/y ), .f(nea) );
    and3_4 \U881/U20/U9  ( .x(nca), .a(\U881/nack[1] ), .b(\U881/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U881/U18/U5  ( .x(\U881/nack[0] ), .a(\cl[3] ), .b(\cl[0] ) );
    nor2_1 \U881/U19/U5  ( .x(\U881/nack[1] ), .a(\cl[1] ), .b(\cl[2] ) );
    ao222_2 \U881/U15_0_/U19/U1/U1  ( .x(\cl[0] ), .a(\c[0] ), .b(ncla), .c(
        \c[0] ), .d(\cl[0] ), .e(ncla), .f(\cl[0] ) );
    ao222_2 \U881/U15_1_/U19/U1/U1  ( .x(\cl[1] ), .a(\c[1] ), .b(ncla), .c(
        \c[1] ), .d(\cl[1] ), .e(ncla), .f(\cl[1] ) );
    ao222_2 \U881/U15_2_/U19/U1/U1  ( .x(\cl[2] ), .a(\c[2] ), .b(ncla), .c(
        \c[2] ), .d(\cl[2] ), .e(ncla), .f(\cl[2] ) );
    ao222_2 \U881/U15_3_/U19/U1/U1  ( .x(\cl[3] ), .a(\c[3] ), .b(ncla), .c(
        \c[3] ), .d(\cl[3] ), .e(ncla), .f(\cl[3] ) );
    and2_5 U1 ( .x(n1), .a(nbReset), .b(noa) );
    and2_3 U2 ( .x(net135), .a(nbReset), .b(noa) );
endmodule


module chain_dr2fr_byte_2 ( eop_ack, ia, o, eop, ih, il, nReset, noa );
output [4:0] o;
input  [7:0] ih;
input  [7:0] il;
input  eop, nReset, noa;
output eop_ack, ia;
    wire eop_pass, nhighack, nlowack, \twobitack[2] , \twobitack[3] , 
        \twobitack[0] , \twobitack[1] , xsel, ysel, nxa, nyla, nbReset, nya, 
        \y[3] , \y[2] , \y[1] , \y[0] , \yl[3] , \yl[2] , \yl[1] , \yl[0] , 
        \cdh[0] , \cdh[1] , \cdl[0] , \cdl[1] , net193, \cdh[2] , \cdh[3] , 
        \cdl[2] , \cdl[3] , net195, bsel, dsel, nba, bg, nda, dg, asel, csel, 
        naa, ag, nca, cg, \d[3] , \d[2] , \d[1] , \d[0] , \b[3] , \b[2] , 
        \b[1] , \b[0] , \x[3] , \x[2] , \x[1] , \x[0] , \c[3] , \c[2] , \c[1] , 
        \c[0] , \a[3] , \a[2] , \a[1] , \a[0] , net194, net199, \U1018/Z , 
        \U1270/net190 , \U1270/net191 , \U1270/net192 , \U1270/net189 , 
        \U1270/U1141/Z , \U1268/net190 , \U1268/net191 , \U1268/net192 , 
        \U1268/net189 , \U1268/U1141/Z , \U1224/nack[0] , \U1224/nack[1] , 
        \U1224/net4 , \U1224/U1125/U28/U1/clr , \U1224/U1125/U28/U1/set , 
        \U1224/U1122/U28/U1/clr , \U1224/U1122/U28/U1/set , 
        \U1224/U916_0_/U25/U1/clr , \U1224/U916_0_/U25/U1/ob , 
        \U1224/U916_1_/U25/U1/clr , \U1224/U916_1_/U25/U1/ob , 
        \U1224/U916_2_/U25/U1/clr , \U1224/U916_2_/U25/U1/ob , 
        \U1224/U916_3_/U25/U1/clr , \U1224/U916_3_/U25/U1/ob , \U1209/nack[0] , 
        \U1209/nack[1] , \U1209/net4 , \U1209/U1125/U28/U1/clr , 
        \U1209/U1125/U28/U1/set , \U1209/U1122/U28/U1/clr , 
        \U1209/U1122/U28/U1/set , \U1209/U916_0_/U25/U1/clr , 
        \U1209/U916_0_/U25/U1/ob , \U1209/U916_1_/U25/U1/clr , 
        \U1209/U916_1_/U25/U1/ob , \U1209/U916_2_/U25/U1/clr , 
        \U1209/U916_2_/U25/U1/ob , \U1209/U916_3_/U25/U1/clr , 
        \U1209/U916_3_/U25/U1/ob , \U1213/nack[0] , \U1213/nack[1] , 
        \U1213/net4 , \U1213/U1125/U28/U1/clr , \U1213/U1125/U28/U1/set , 
        \U1213/U1122/U28/U1/clr , \U1213/U1122/U28/U1/set , 
        \U1213/U916_0_/U25/U1/clr , \U1213/U916_0_/U25/U1/ob , 
        \U1213/U916_1_/U25/U1/clr , \U1213/U916_1_/U25/U1/ob , 
        \U1213/U916_2_/U25/U1/clr , \U1213/U916_2_/U25/U1/ob , 
        \U1213/U916_3_/U25/U1/clr , \U1213/U916_3_/U25/U1/ob , \U1296/ng , 
        \U1296/U1384/Z , \U1296/U1386/U25/U1/clr , \U1296/U1386/U25/U1/ob , 
        \U1298/ng , \U1298/U1384/Z , \U1298/U1386/U25/U1/clr , 
        \U1298/U1386/U25/U1/ob , \U1306/ng , \U1306/U1384/Z , 
        \U1306/U1386/U25/U1/clr , \U1306/U1386/U25/U1/ob , \U1295/ng , 
        \U1295/U1384/Z , \U1295/U1386/U25/U1/clr , \U1295/U1386/U25/U1/ob , 
        \U1297/s , \U1297/nback , \U1297/r , \U1297/naack , \U1297/reset , 
        \U1297/U1128/U28/U1/clr , \U1297/U1128/U28/U1/set , 
        \U1297/U1127/U28/U1/clr , \U1297/U1127/U28/U1/set , \U1300/s , 
        \U1300/nback , \U1300/r , \U1300/naack , \U1300/reset , 
        \U1300/U1128/U28/U1/clr , \U1300/U1128/U28/U1/set , 
        \U1300/U1127/U28/U1/clr , \U1300/U1127/U28/U1/set , \U1289/bnreset , 
        \U1289/U1150/U28/U1/clr , \U1289/U1150/U28/U1/set , 
        \U1289/U1152/U28/U1/clr , \U1289/U1152/U28/U1/set , 
        \U1289/U1149/U28/U1/clr , \U1289/U1149/U28/U1/set , 
        \U1289/U1151/U28/U1/clr , \U1289/U1151/U28/U1/set , 
        \U1289/U1148/net190 , \U1289/U1148/net191 , \U1289/U1148/net192 , 
        \U1289/U1148/net189 , \U1289/U1148/U1141/Z , \U1271/bnreset , 
        \U1271/U1150/U28/U1/clr , \U1271/U1150/U28/U1/set , 
        \U1271/U1152/U28/U1/clr , \U1271/U1152/U28/U1/set , 
        \U1271/U1149/U28/U1/clr , \U1271/U1149/U28/U1/set , 
        \U1271/U1151/U28/U1/clr , \U1271/U1151/U28/U1/set , 
        \U1271/U1148/net190 , \U1271/U1148/net191 , \U1271/U1148/net192 , 
        \U1271/U1148/net189 , \U1271/U1148/U1141/Z , \U1225/naack , \U1225/r , 
        \U1225/s , \U1225/nback , \U1225/reset , \U1308/nack[1] , 
        \U1308/nack[0] ;
    assign o[4] = eop_ack;
    buf_2 U1231 ( .x(nbReset), .a(nReset) );
    and3_1 \U1194/U9  ( .x(eop_pass), .a(nxa), .b(naa), .c(eop) );
    ao222_1 \U1301/U18/U1/U1  ( .x(nlowack), .a(\twobitack[0] ), .b(
        \twobitack[1] ), .c(\twobitack[0] ), .d(nlowack), .e(\twobitack[1] ), 
        .f(nlowack) );
    ao222_1 \U1302/U18/U1/U1  ( .x(nhighack), .a(\twobitack[2] ), .b(
        \twobitack[3] ), .c(\twobitack[2] ), .d(nhighack), .e(\twobitack[3] ), 
        .f(nhighack) );
    aoi222_1 \U1018/U30/U1  ( .x(ia), .a(nhighack), .b(nlowack), .c(nhighack), 
        .d(\U1018/Z ), .e(nlowack), .f(\U1018/Z ) );
    inv_1 \U1018/U30/Uinv  ( .x(\U1018/Z ), .a(ia) );
    ao222_2 \U1038/U19/U1/U1  ( .x(eop_ack), .a(eop_pass), .b(noa), .c(
        eop_pass), .d(eop_ack), .e(noa), .f(eop_ack) );
    inv_1 \U1270/U1147/U3  ( .x(\U1270/net189 ), .a(nbReset) );
    nor2_1 \U1270/U582/U5  ( .x(\U1270/net192 ), .a(il[4]), .b(ih[4]) );
    nor2_1 \U1270/U580/U5  ( .x(\U1270/net191 ), .a(il[5]), .b(ih[5]) );
    nor2_2 \U1270/U1146/U6  ( .x(net199), .a(\U1270/net190 ), .b(
        \U1270/net189 ) );
    aoi222_1 \U1270/U1141/U30/U1  ( .x(\U1270/net190 ), .a(\U1270/net191 ), 
        .b(\U1270/net192 ), .c(\U1270/net191 ), .d(\U1270/U1141/Z ), .e(
        \U1270/net192 ), .f(\U1270/U1141/Z ) );
    inv_1 \U1270/U1141/U30/Uinv  ( .x(\U1270/U1141/Z ), .a(\U1270/net190 ) );
    inv_1 \U1268/U1147/U3  ( .x(\U1268/net189 ), .a(nbReset) );
    nor2_1 \U1268/U582/U5  ( .x(\U1268/net192 ), .a(il[6]), .b(ih[6]) );
    nor2_1 \U1268/U580/U5  ( .x(\U1268/net191 ), .a(il[7]), .b(ih[7]) );
    nor2_2 \U1268/U1146/U6  ( .x(net194), .a(\U1268/net190 ), .b(
        \U1268/net189 ) );
    aoi222_1 \U1268/U1141/U30/U1  ( .x(\U1268/net190 ), .a(\U1268/net191 ), 
        .b(\U1268/net192 ), .c(\U1268/net191 ), .d(\U1268/U1141/Z ), .e(
        \U1268/net192 ), .f(\U1268/U1141/Z ) );
    inv_1 \U1268/U1141/U30/Uinv  ( .x(\U1268/U1141/Z ), .a(\U1268/net190 ) );
    nor2_1 \U1224/U1128/U5  ( .x(\U1224/nack[0] ), .a(\x[3] ), .b(\x[2] ) );
    nor3_1 \U1224/U1127/U7  ( .x(\U1224/nack[1] ), .a(\x[1] ), .b(\U1224/net4 
        ), .c(\x[0] ) );
    inv_1 \U1224/U907/U3  ( .x(\U1224/net4 ), .a(nbReset) );
    aoai211_1 \U1224/U1125/U28/U1/U1  ( .x(\U1224/U1125/U28/U1/clr ), .a(
        \U1224/nack[1] ), .b(\U1224/nack[0] ), .c(asel), .d(naa) );
    nand3_1 \U1224/U1125/U28/U1/U2  ( .x(\U1224/U1125/U28/U1/set ), .a(asel), 
        .b(\U1224/nack[1] ), .c(\U1224/nack[0] ) );
    nand2_2 \U1224/U1125/U28/U1/U3  ( .x(naa), .a(\U1224/U1125/U28/U1/clr ), 
        .b(\U1224/U1125/U28/U1/set ) );
    aoai211_1 \U1224/U1122/U28/U1/U1  ( .x(\U1224/U1122/U28/U1/clr ), .a(
        \U1224/nack[0] ), .b(\U1224/nack[1] ), .c(csel), .d(nca) );
    nand3_1 \U1224/U1122/U28/U1/U2  ( .x(\U1224/U1122/U28/U1/set ), .a(csel), 
        .b(\U1224/nack[0] ), .c(\U1224/nack[1] ) );
    nand2_2 \U1224/U1122/U28/U1/U3  ( .x(nca), .a(\U1224/U1122/U28/U1/clr ), 
        .b(\U1224/U1122/U28/U1/set ) );
    oa31_1 \U1224/U916_0_/U25/U1/Uclr  ( .x(\U1224/U916_0_/U25/U1/clr ), .a(
        nxa), .b(\a[0] ), .c(\c[0] ), .d(\x[0] ) );
    oaoi211_1 \U1224/U916_0_/U25/U1/Uaoi  ( .x(\U1224/U916_0_/U25/U1/ob ), .a(
        \a[0] ), .b(\c[0] ), .c(nxa), .d(\U1224/U916_0_/U25/U1/clr ) );
    inv_2 \U1224/U916_0_/U25/U1/Ui  ( .x(\x[0] ), .a(\U1224/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_1_/U25/U1/Uclr  ( .x(\U1224/U916_1_/U25/U1/clr ), .a(
        nxa), .b(\a[1] ), .c(\c[1] ), .d(\x[1] ) );
    oaoi211_1 \U1224/U916_1_/U25/U1/Uaoi  ( .x(\U1224/U916_1_/U25/U1/ob ), .a(
        \a[1] ), .b(\c[1] ), .c(nxa), .d(\U1224/U916_1_/U25/U1/clr ) );
    inv_2 \U1224/U916_1_/U25/U1/Ui  ( .x(\x[1] ), .a(\U1224/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_2_/U25/U1/Uclr  ( .x(\U1224/U916_2_/U25/U1/clr ), .a(
        nxa), .b(\a[2] ), .c(\c[2] ), .d(\x[2] ) );
    oaoi211_1 \U1224/U916_2_/U25/U1/Uaoi  ( .x(\U1224/U916_2_/U25/U1/ob ), .a(
        \a[2] ), .b(\c[2] ), .c(nxa), .d(\U1224/U916_2_/U25/U1/clr ) );
    inv_2 \U1224/U916_2_/U25/U1/Ui  ( .x(\x[2] ), .a(\U1224/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_3_/U25/U1/Uclr  ( .x(\U1224/U916_3_/U25/U1/clr ), .a(
        nxa), .b(\a[3] ), .c(\c[3] ), .d(\x[3] ) );
    oaoi211_1 \U1224/U916_3_/U25/U1/Uaoi  ( .x(\U1224/U916_3_/U25/U1/ob ), .a(
        \a[3] ), .b(\c[3] ), .c(nxa), .d(\U1224/U916_3_/U25/U1/clr ) );
    inv_2 \U1224/U916_3_/U25/U1/Ui  ( .x(\x[3] ), .a(\U1224/U916_3_/U25/U1/ob 
        ) );
    nor2_1 \U1209/U1128/U5  ( .x(\U1209/nack[0] ), .a(o[3]), .b(o[2]) );
    nor3_1 \U1209/U1127/U7  ( .x(\U1209/nack[1] ), .a(o[1]), .b(\U1209/net4 ), 
        .c(o[0]) );
    inv_1 \U1209/U907/U3  ( .x(\U1209/net4 ), .a(nbReset) );
    aoai211_1 \U1209/U1125/U28/U1/U1  ( .x(\U1209/U1125/U28/U1/clr ), .a(
        \U1209/nack[1] ), .b(\U1209/nack[0] ), .c(xsel), .d(nxa) );
    nand3_1 \U1209/U1125/U28/U1/U2  ( .x(\U1209/U1125/U28/U1/set ), .a(xsel), 
        .b(\U1209/nack[1] ), .c(\U1209/nack[0] ) );
    nand2_2 \U1209/U1125/U28/U1/U3  ( .x(nxa), .a(\U1209/U1125/U28/U1/clr ), 
        .b(\U1209/U1125/U28/U1/set ) );
    aoai211_1 \U1209/U1122/U28/U1/U1  ( .x(\U1209/U1122/U28/U1/clr ), .a(
        \U1209/nack[0] ), .b(\U1209/nack[1] ), .c(ysel), .d(nyla) );
    nand3_1 \U1209/U1122/U28/U1/U2  ( .x(\U1209/U1122/U28/U1/set ), .a(ysel), 
        .b(\U1209/nack[0] ), .c(\U1209/nack[1] ) );
    nand2_2 \U1209/U1122/U28/U1/U3  ( .x(nyla), .a(\U1209/U1122/U28/U1/clr ), 
        .b(\U1209/U1122/U28/U1/set ) );
    oa31_1 \U1209/U916_0_/U25/U1/Uclr  ( .x(\U1209/U916_0_/U25/U1/clr ), .a(
        noa), .b(\x[0] ), .c(\yl[0] ), .d(o[0]) );
    oaoi211_1 \U1209/U916_0_/U25/U1/Uaoi  ( .x(\U1209/U916_0_/U25/U1/ob ), .a(
        \x[0] ), .b(\yl[0] ), .c(noa), .d(\U1209/U916_0_/U25/U1/clr ) );
    inv_2 \U1209/U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U1209/U916_0_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_1_/U25/U1/Uclr  ( .x(\U1209/U916_1_/U25/U1/clr ), .a(
        noa), .b(\x[1] ), .c(\yl[1] ), .d(o[1]) );
    oaoi211_1 \U1209/U916_1_/U25/U1/Uaoi  ( .x(\U1209/U916_1_/U25/U1/ob ), .a(
        \x[1] ), .b(\yl[1] ), .c(noa), .d(\U1209/U916_1_/U25/U1/clr ) );
    inv_2 \U1209/U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U1209/U916_1_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_2_/U25/U1/Uclr  ( .x(\U1209/U916_2_/U25/U1/clr ), .a(
        noa), .b(\x[2] ), .c(\yl[2] ), .d(o[2]) );
    oaoi211_1 \U1209/U916_2_/U25/U1/Uaoi  ( .x(\U1209/U916_2_/U25/U1/ob ), .a(
        \x[2] ), .b(\yl[2] ), .c(noa), .d(\U1209/U916_2_/U25/U1/clr ) );
    inv_2 \U1209/U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U1209/U916_2_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_3_/U25/U1/Uclr  ( .x(\U1209/U916_3_/U25/U1/clr ), .a(
        noa), .b(\x[3] ), .c(\yl[3] ), .d(o[3]) );
    oaoi211_1 \U1209/U916_3_/U25/U1/Uaoi  ( .x(\U1209/U916_3_/U25/U1/ob ), .a(
        \x[3] ), .b(\yl[3] ), .c(noa), .d(\U1209/U916_3_/U25/U1/clr ) );
    inv_2 \U1209/U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U1209/U916_3_/U25/U1/ob )
         );
    nor2_1 \U1213/U1128/U5  ( .x(\U1213/nack[0] ), .a(\y[3] ), .b(\y[2] ) );
    nor3_1 \U1213/U1127/U7  ( .x(\U1213/nack[1] ), .a(\y[1] ), .b(\U1213/net4 
        ), .c(\y[0] ) );
    inv_1 \U1213/U907/U3  ( .x(\U1213/net4 ), .a(nbReset) );
    aoai211_1 \U1213/U1125/U28/U1/U1  ( .x(\U1213/U1125/U28/U1/clr ), .a(
        \U1213/nack[1] ), .b(\U1213/nack[0] ), .c(bsel), .d(nba) );
    nand3_1 \U1213/U1125/U28/U1/U2  ( .x(\U1213/U1125/U28/U1/set ), .a(bsel), 
        .b(\U1213/nack[1] ), .c(\U1213/nack[0] ) );
    nand2_2 \U1213/U1125/U28/U1/U3  ( .x(nba), .a(\U1213/U1125/U28/U1/clr ), 
        .b(\U1213/U1125/U28/U1/set ) );
    aoai211_1 \U1213/U1122/U28/U1/U1  ( .x(\U1213/U1122/U28/U1/clr ), .a(
        \U1213/nack[0] ), .b(\U1213/nack[1] ), .c(dsel), .d(nda) );
    nand3_1 \U1213/U1122/U28/U1/U2  ( .x(\U1213/U1122/U28/U1/set ), .a(dsel), 
        .b(\U1213/nack[0] ), .c(\U1213/nack[1] ) );
    nand2_2 \U1213/U1122/U28/U1/U3  ( .x(nda), .a(\U1213/U1122/U28/U1/clr ), 
        .b(\U1213/U1122/U28/U1/set ) );
    oa31_1 \U1213/U916_0_/U25/U1/Uclr  ( .x(\U1213/U916_0_/U25/U1/clr ), .a(
        nya), .b(\b[0] ), .c(\d[0] ), .d(\y[0] ) );
    oaoi211_1 \U1213/U916_0_/U25/U1/Uaoi  ( .x(\U1213/U916_0_/U25/U1/ob ), .a(
        \b[0] ), .b(\d[0] ), .c(nya), .d(\U1213/U916_0_/U25/U1/clr ) );
    inv_2 \U1213/U916_0_/U25/U1/Ui  ( .x(\y[0] ), .a(\U1213/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_1_/U25/U1/Uclr  ( .x(\U1213/U916_1_/U25/U1/clr ), .a(
        nya), .b(\b[1] ), .c(\d[1] ), .d(\y[1] ) );
    oaoi211_1 \U1213/U916_1_/U25/U1/Uaoi  ( .x(\U1213/U916_1_/U25/U1/ob ), .a(
        \b[1] ), .b(\d[1] ), .c(nya), .d(\U1213/U916_1_/U25/U1/clr ) );
    inv_2 \U1213/U916_1_/U25/U1/Ui  ( .x(\y[1] ), .a(\U1213/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_2_/U25/U1/Uclr  ( .x(\U1213/U916_2_/U25/U1/clr ), .a(
        nya), .b(\b[2] ), .c(\d[2] ), .d(\y[2] ) );
    oaoi211_1 \U1213/U916_2_/U25/U1/Uaoi  ( .x(\U1213/U916_2_/U25/U1/ob ), .a(
        \b[2] ), .b(\d[2] ), .c(nya), .d(\U1213/U916_2_/U25/U1/clr ) );
    inv_2 \U1213/U916_2_/U25/U1/Ui  ( .x(\y[2] ), .a(\U1213/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_3_/U25/U1/Uclr  ( .x(\U1213/U916_3_/U25/U1/clr ), .a(
        nya), .b(\b[3] ), .c(\d[3] ), .d(\y[3] ) );
    oaoi211_1 \U1213/U916_3_/U25/U1/Uaoi  ( .x(\U1213/U916_3_/U25/U1/ob ), .a(
        \b[3] ), .b(\d[3] ), .c(nya), .d(\U1213/U916_3_/U25/U1/clr ) );
    inv_2 \U1213/U916_3_/U25/U1/Ui  ( .x(\y[3] ), .a(\U1213/U916_3_/U25/U1/ob 
        ) );
    and3_2 \U1210/U1138/U9  ( .x(\d[3] ), .a(\cdh[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1137/U9  ( .x(\d[2] ), .a(\cdl[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1139/U9  ( .x(\d[1] ), .a(\cdh[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1210/U1136/U9  ( .x(\d[0] ), .a(\cdl[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1162/U1138/U9  ( .x(\a[3] ), .a(ih[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1137/U9  ( .x(\a[2] ), .a(il[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1139/U9  ( .x(\a[1] ), .a(ih[6]), .b(naa), .c(il[7]) );
    and3_2 \U1162/U1136/U9  ( .x(\a[0] ), .a(il[6]), .b(naa), .c(il[7]) );
    and3_2 \U1211/U1138/U9  ( .x(\b[3] ), .a(ih[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1137/U9  ( .x(\b[2] ), .a(il[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1139/U9  ( .x(\b[1] ), .a(ih[4]), .b(nba), .c(il[5]) );
    and3_2 \U1211/U1136/U9  ( .x(\b[0] ), .a(il[4]), .b(nba), .c(il[5]) );
    and3_2 \U1163/U1138/U9  ( .x(\c[3] ), .a(\cdh[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1137/U9  ( .x(\c[2] ), .a(\cdl[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1139/U9  ( .x(\c[1] ), .a(\cdh[2] ), .b(nca), .c(\cdl[3] )
         );
    and3_2 \U1163/U1136/U9  ( .x(\c[0] ), .a(\cdl[2] ), .b(nca), .c(\cdl[3] )
         );
    and2_1 \U1296/U1385/U8  ( .x(cg), .a(nbReset), .b(\U1296/ng ) );
    aoi222_1 \U1296/U1384/U30/U1  ( .x(\U1296/ng ), .a(nca), .b(net195), .c(
        nca), .d(\U1296/U1384/Z ), .e(net195), .f(\U1296/U1384/Z ) );
    inv_1 \U1296/U1384/U30/Uinv  ( .x(\U1296/U1384/Z ), .a(\U1296/ng ) );
    oa31_1 \U1296/U1386/U25/U1/Uclr  ( .x(\U1296/U1386/U25/U1/clr ), .a(
        \twobitack[2] ), .b(cg), .c(nca), .d(net195) );
    oaoi211_1 \U1296/U1386/U25/U1/Uaoi  ( .x(\U1296/U1386/U25/U1/ob ), .a(cg), 
        .b(nca), .c(\twobitack[2] ), .d(\U1296/U1386/U25/U1/clr ) );
    inv_2 \U1296/U1386/U25/U1/Ui  ( .x(net195), .a(\U1296/U1386/U25/U1/ob ) );
    and2_1 \U1298/U1385/U8  ( .x(dg), .a(nbReset), .b(\U1298/ng ) );
    aoi222_1 \U1298/U1384/U30/U1  ( .x(\U1298/ng ), .a(nda), .b(net193), .c(
        nda), .d(\U1298/U1384/Z ), .e(net193), .f(\U1298/U1384/Z ) );
    inv_1 \U1298/U1384/U30/Uinv  ( .x(\U1298/U1384/Z ), .a(\U1298/ng ) );
    oa31_1 \U1298/U1386/U25/U1/Uclr  ( .x(\U1298/U1386/U25/U1/clr ), .a(
        \twobitack[0] ), .b(dg), .c(nda), .d(net193) );
    oaoi211_1 \U1298/U1386/U25/U1/Uaoi  ( .x(\U1298/U1386/U25/U1/ob ), .a(dg), 
        .b(nda), .c(\twobitack[0] ), .d(\U1298/U1386/U25/U1/clr ) );
    inv_2 \U1298/U1386/U25/U1/Ui  ( .x(net193), .a(\U1298/U1386/U25/U1/ob ) );
    and2_1 \U1306/U1385/U8  ( .x(bg), .a(nbReset), .b(\U1306/ng ) );
    aoi222_1 \U1306/U1384/U30/U1  ( .x(\U1306/ng ), .a(nba), .b(\twobitack[1] 
        ), .c(nba), .d(\U1306/U1384/Z ), .e(\twobitack[1] ), .f(
        \U1306/U1384/Z ) );
    inv_1 \U1306/U1384/U30/Uinv  ( .x(\U1306/U1384/Z ), .a(\U1306/ng ) );
    oa31_1 \U1306/U1386/U25/U1/Uclr  ( .x(\U1306/U1386/U25/U1/clr ), .a(net199
        ), .b(bg), .c(nba), .d(\twobitack[1] ) );
    oaoi211_1 \U1306/U1386/U25/U1/Uaoi  ( .x(\U1306/U1386/U25/U1/ob ), .a(bg), 
        .b(nba), .c(net199), .d(\U1306/U1386/U25/U1/clr ) );
    inv_2 \U1306/U1386/U25/U1/Ui  ( .x(\twobitack[1] ), .a(
        \U1306/U1386/U25/U1/ob ) );
    and2_1 \U1295/U1385/U8  ( .x(ag), .a(nbReset), .b(\U1295/ng ) );
    aoi222_1 \U1295/U1384/U30/U1  ( .x(\U1295/ng ), .a(naa), .b(\twobitack[3] 
        ), .c(naa), .d(\U1295/U1384/Z ), .e(\twobitack[3] ), .f(
        \U1295/U1384/Z ) );
    inv_1 \U1295/U1384/U30/Uinv  ( .x(\U1295/U1384/Z ), .a(\U1295/ng ) );
    oa31_1 \U1295/U1386/U25/U1/Uclr  ( .x(\U1295/U1386/U25/U1/clr ), .a(net194
        ), .b(ag), .c(naa), .d(\twobitack[3] ) );
    oaoi211_1 \U1295/U1386/U25/U1/Uaoi  ( .x(\U1295/U1386/U25/U1/ob ), .a(ag), 
        .b(naa), .c(net194), .d(\U1295/U1386/U25/U1/clr ) );
    inv_2 \U1295/U1386/U25/U1/Ui  ( .x(\twobitack[3] ), .a(
        \U1295/U1386/U25/U1/ob ) );
    nand2_1 \U1297/U1131/U5  ( .x(\U1297/s ), .a(\U1297/r ), .b(\U1297/nback )
         );
    nand2_1 \U1297/U1103/U5  ( .x(\U1297/r ), .a(\U1297/naack ), .b(\U1297/s )
         );
    inv_1 \U1297/U1111/U3  ( .x(\U1297/reset ), .a(nbReset) );
    inv_1 \U1297/U1112/U3  ( .x(\U1297/naack ), .a(naa) );
    nor2_1 \U1297/U1130/U5  ( .x(\U1297/nback ), .a(nca), .b(\U1297/reset ) );
    aoai211_1 \U1297/U1128/U28/U1/U1  ( .x(\U1297/U1128/U28/U1/clr ), .a(
        \U1297/r ), .b(\U1297/naack ), .c(cg), .d(csel) );
    nand3_1 \U1297/U1128/U28/U1/U2  ( .x(\U1297/U1128/U28/U1/set ), .a(cg), 
        .b(\U1297/r ), .c(\U1297/naack ) );
    nand2_2 \U1297/U1128/U28/U1/U3  ( .x(csel), .a(\U1297/U1128/U28/U1/clr ), 
        .b(\U1297/U1128/U28/U1/set ) );
    aoai211_1 \U1297/U1127/U28/U1/U1  ( .x(\U1297/U1127/U28/U1/clr ), .a(
        \U1297/s ), .b(\U1297/nback ), .c(ag), .d(asel) );
    nand3_1 \U1297/U1127/U28/U1/U2  ( .x(\U1297/U1127/U28/U1/set ), .a(ag), 
        .b(\U1297/s ), .c(\U1297/nback ) );
    nand2_2 \U1297/U1127/U28/U1/U3  ( .x(asel), .a(\U1297/U1127/U28/U1/clr ), 
        .b(\U1297/U1127/U28/U1/set ) );
    nand2_1 \U1300/U1131/U5  ( .x(\U1300/s ), .a(\U1300/r ), .b(\U1300/nback )
         );
    nand2_1 \U1300/U1103/U5  ( .x(\U1300/r ), .a(\U1300/naack ), .b(\U1300/s )
         );
    inv_1 \U1300/U1111/U3  ( .x(\U1300/reset ), .a(nbReset) );
    inv_1 \U1300/U1112/U3  ( .x(\U1300/naack ), .a(nba) );
    nor2_1 \U1300/U1130/U5  ( .x(\U1300/nback ), .a(nda), .b(\U1300/reset ) );
    aoai211_1 \U1300/U1128/U28/U1/U1  ( .x(\U1300/U1128/U28/U1/clr ), .a(
        \U1300/r ), .b(\U1300/naack ), .c(dg), .d(dsel) );
    nand3_1 \U1300/U1128/U28/U1/U2  ( .x(\U1300/U1128/U28/U1/set ), .a(dg), 
        .b(\U1300/r ), .c(\U1300/naack ) );
    nand2_2 \U1300/U1128/U28/U1/U3  ( .x(dsel), .a(\U1300/U1128/U28/U1/clr ), 
        .b(\U1300/U1128/U28/U1/set ) );
    aoai211_1 \U1300/U1127/U28/U1/U1  ( .x(\U1300/U1127/U28/U1/clr ), .a(
        \U1300/s ), .b(\U1300/nback ), .c(bg), .d(bsel) );
    nand3_1 \U1300/U1127/U28/U1/U2  ( .x(\U1300/U1127/U28/U1/set ), .a(bg), 
        .b(\U1300/s ), .c(\U1300/nback ) );
    nand2_2 \U1300/U1127/U28/U1/U3  ( .x(bsel), .a(\U1300/U1127/U28/U1/clr ), 
        .b(\U1300/U1127/U28/U1/set ) );
    aoai211_1 \U1289/U1150/U28/U1/U1  ( .x(\U1289/U1150/U28/U1/clr ), .a(il[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[2] ) );
    nand3_1 \U1289/U1150/U28/U1/U2  ( .x(\U1289/U1150/U28/U1/set ), .a(net195), 
        .b(il[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1150/U28/U1/U3  ( .x(\cdl[2] ), .a(
        \U1289/U1150/U28/U1/clr ), .b(\U1289/U1150/U28/U1/set ) );
    aoai211_1 \U1289/U1152/U28/U1/U1  ( .x(\U1289/U1152/U28/U1/clr ), .a(il[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[3] ) );
    nand3_1 \U1289/U1152/U28/U1/U2  ( .x(\U1289/U1152/U28/U1/set ), .a(net195), 
        .b(il[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1152/U28/U1/U3  ( .x(\cdl[3] ), .a(
        \U1289/U1152/U28/U1/clr ), .b(\U1289/U1152/U28/U1/set ) );
    aoai211_1 \U1289/U1149/U28/U1/U1  ( .x(\U1289/U1149/U28/U1/clr ), .a(ih[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[2] ) );
    nand3_1 \U1289/U1149/U28/U1/U2  ( .x(\U1289/U1149/U28/U1/set ), .a(net195), 
        .b(ih[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1149/U28/U1/U3  ( .x(\cdh[2] ), .a(
        \U1289/U1149/U28/U1/clr ), .b(\U1289/U1149/U28/U1/set ) );
    aoai211_1 \U1289/U1151/U28/U1/U1  ( .x(\U1289/U1151/U28/U1/clr ), .a(ih[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[3] ) );
    nand3_1 \U1289/U1151/U28/U1/U2  ( .x(\U1289/U1151/U28/U1/set ), .a(net195), 
        .b(ih[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1151/U28/U1/U3  ( .x(\cdh[3] ), .a(
        \U1289/U1151/U28/U1/clr ), .b(\U1289/U1151/U28/U1/set ) );
    inv_1 \U1289/U1148/U1147/U3  ( .x(\U1289/U1148/net189 ), .a(
        \U1289/bnreset ) );
    nor2_1 \U1289/U1148/U582/U5  ( .x(\U1289/U1148/net192 ), .a(\cdl[3] ), .b(
        \cdh[3] ) );
    nor2_1 \U1289/U1148/U580/U5  ( .x(\U1289/U1148/net191 ), .a(\cdl[2] ), .b(
        \cdh[2] ) );
    nor2_2 \U1289/U1148/U1146/U6  ( .x(\twobitack[2] ), .a(
        \U1289/U1148/net190 ), .b(\U1289/U1148/net189 ) );
    aoi222_1 \U1289/U1148/U1141/U30/U1  ( .x(\U1289/U1148/net190 ), .a(
        \U1289/U1148/net191 ), .b(\U1289/U1148/net192 ), .c(
        \U1289/U1148/net191 ), .d(\U1289/U1148/U1141/Z ), .e(
        \U1289/U1148/net192 ), .f(\U1289/U1148/U1141/Z ) );
    inv_1 \U1289/U1148/U1141/U30/Uinv  ( .x(\U1289/U1148/U1141/Z ), .a(
        \U1289/U1148/net190 ) );
    aoai211_1 \U1271/U1150/U28/U1/U1  ( .x(\U1271/U1150/U28/U1/clr ), .a(il[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[0] ) );
    nand3_1 \U1271/U1150/U28/U1/U2  ( .x(\U1271/U1150/U28/U1/set ), .a(net193), 
        .b(il[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1150/U28/U1/U3  ( .x(\cdl[0] ), .a(
        \U1271/U1150/U28/U1/clr ), .b(\U1271/U1150/U28/U1/set ) );
    aoai211_1 \U1271/U1152/U28/U1/U1  ( .x(\U1271/U1152/U28/U1/clr ), .a(il[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[1] ) );
    nand3_1 \U1271/U1152/U28/U1/U2  ( .x(\U1271/U1152/U28/U1/set ), .a(net193), 
        .b(il[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1152/U28/U1/U3  ( .x(\cdl[1] ), .a(
        \U1271/U1152/U28/U1/clr ), .b(\U1271/U1152/U28/U1/set ) );
    aoai211_1 \U1271/U1149/U28/U1/U1  ( .x(\U1271/U1149/U28/U1/clr ), .a(ih[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[0] ) );
    nand3_1 \U1271/U1149/U28/U1/U2  ( .x(\U1271/U1149/U28/U1/set ), .a(net193), 
        .b(ih[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1149/U28/U1/U3  ( .x(\cdh[0] ), .a(
        \U1271/U1149/U28/U1/clr ), .b(\U1271/U1149/U28/U1/set ) );
    aoai211_1 \U1271/U1151/U28/U1/U1  ( .x(\U1271/U1151/U28/U1/clr ), .a(ih[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[1] ) );
    nand3_1 \U1271/U1151/U28/U1/U2  ( .x(\U1271/U1151/U28/U1/set ), .a(net193), 
        .b(ih[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1151/U28/U1/U3  ( .x(\cdh[1] ), .a(
        \U1271/U1151/U28/U1/clr ), .b(\U1271/U1151/U28/U1/set ) );
    inv_1 \U1271/U1148/U1147/U3  ( .x(\U1271/U1148/net189 ), .a(
        \U1271/bnreset ) );
    nor2_1 \U1271/U1148/U582/U5  ( .x(\U1271/U1148/net192 ), .a(\cdl[1] ), .b(
        \cdh[1] ) );
    nor2_1 \U1271/U1148/U580/U5  ( .x(\U1271/U1148/net191 ), .a(\cdl[0] ), .b(
        \cdh[0] ) );
    nor2_2 \U1271/U1148/U1146/U6  ( .x(\twobitack[0] ), .a(
        \U1271/U1148/net190 ), .b(\U1271/U1148/net189 ) );
    aoi222_1 \U1271/U1148/U1141/U30/U1  ( .x(\U1271/U1148/net190 ), .a(
        \U1271/U1148/net191 ), .b(\U1271/U1148/net192 ), .c(
        \U1271/U1148/net191 ), .d(\U1271/U1148/U1141/Z ), .e(
        \U1271/U1148/net192 ), .f(\U1271/U1148/U1141/Z ) );
    inv_1 \U1271/U1148/U1141/U30/Uinv  ( .x(\U1271/U1148/U1141/Z ), .a(
        \U1271/U1148/net190 ) );
    nand2_1 \U1225/U1128/U5  ( .x(\U1225/s ), .a(\U1225/r ), .b(\U1225/nback )
         );
    nand2_1 \U1225/U1103/U5  ( .x(\U1225/r ), .a(\U1225/naack ), .b(\U1225/s )
         );
    inv_1 \U1225/U1111/U3  ( .x(\U1225/reset ), .a(nbReset) );
    inv_1 \U1225/U1112/U3  ( .x(\U1225/naack ), .a(nxa) );
    nor2_1 \U1225/U1127/U5  ( .x(\U1225/nback ), .a(nyla), .b(\U1225/reset )
         );
    and2_2 \U1225/U1129/U8  ( .x(xsel), .a(\U1225/nback ), .b(\U1225/s ) );
    and2_2 \U1225/U1124/U8  ( .x(ysel), .a(\U1225/r ), .b(\U1225/naack ) );
    and3_4 \U1308/U20/U9  ( .x(nya), .a(\U1308/nack[1] ), .b(\U1308/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U1308/U18/U5  ( .x(\U1308/nack[0] ), .a(\yl[3] ), .b(\yl[0] ) );
    nor2_1 \U1308/U19/U5  ( .x(\U1308/nack[1] ), .a(\yl[1] ), .b(\yl[2] ) );
    ao222_2 \U1308/U15_0_/U19/U1/U1  ( .x(\yl[0] ), .a(\y[0] ), .b(nyla), .c(
        \y[0] ), .d(\yl[0] ), .e(nyla), .f(\yl[0] ) );
    ao222_2 \U1308/U15_1_/U19/U1/U1  ( .x(\yl[1] ), .a(\y[1] ), .b(nyla), .c(
        \y[1] ), .d(\yl[1] ), .e(nyla), .f(\yl[1] ) );
    ao222_2 \U1308/U15_2_/U19/U1/U1  ( .x(\yl[2] ), .a(\y[2] ), .b(nyla), .c(
        \y[2] ), .d(\yl[2] ), .e(nyla), .f(\yl[2] ) );
    ao222_2 \U1308/U15_3_/U19/U1/U1  ( .x(\yl[3] ), .a(\y[3] ), .b(nyla), .c(
        \y[3] ), .d(\yl[3] ), .e(nyla), .f(\yl[3] ) );
    buf_3 U1 ( .x(\U1289/bnreset ), .a(nbReset) );
    buf_3 U2 ( .x(\U1271/bnreset ), .a(nbReset) );
endmodule


module chain_mergepackets_2 ( naa, nba, o, a, b, nReset, noa );
output [4:0] o;
input  [4:0] a;
input  [4:0] b;
input  nReset, noa;
output naa, nba;
    wire \noack[1] , \noack[0] , reset, bsel, as, setb, asel, seta, 
        \U916_0_/U25/U1/clr , \U916_0_/U25/U1/ob , \U916_1_/U25/U1/clr , 
        \U916_1_/U25/U1/ob , \U916_2_/U25/U1/clr , \U916_2_/U25/U1/ob , 
        \U916_3_/U25/U1/clr , \U916_3_/U25/U1/ob ;
    and2_1 \U1155/U8  ( .x(as), .a(seta), .b(asel) );
    nand2_1 \U1145/U5  ( .x(asel), .a(bsel), .b(seta) );
    nand2_1 \U1103/U5  ( .x(bsel), .a(setb), .b(asel) );
    inv_1 \U1135/U3  ( .x(reset), .a(nReset) );
    inv_1 \U1134/U3  ( .x(setb), .a(a[4]) );
    and3_2 \U1154/U9  ( .x(naa), .a(\noack[1] ), .b(\noack[0] ), .c(as) );
    nor3_1 \U1127/U7  ( .x(\noack[0] ), .a(o[1]), .b(reset), .c(o[0]) );
    nor2_1 \U1132/U5  ( .x(\noack[1] ), .a(o[3]), .b(o[2]) );
    oa31_1 \U916_0_/U25/U1/Uclr  ( .x(\U916_0_/U25/U1/clr ), .a(noa), .b(a[0]), 
        .c(b[0]), .d(o[0]) );
    oaoi211_1 \U916_0_/U25/U1/Uaoi  ( .x(\U916_0_/U25/U1/ob ), .a(a[0]), .b(b
        [0]), .c(noa), .d(\U916_0_/U25/U1/clr ) );
    inv_2 \U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U916_0_/U25/U1/ob ) );
    oa31_1 \U916_1_/U25/U1/Uclr  ( .x(\U916_1_/U25/U1/clr ), .a(noa), .b(a[1]), 
        .c(b[1]), .d(o[1]) );
    oaoi211_1 \U916_1_/U25/U1/Uaoi  ( .x(\U916_1_/U25/U1/ob ), .a(a[1]), .b(b
        [1]), .c(noa), .d(\U916_1_/U25/U1/clr ) );
    inv_2 \U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U916_1_/U25/U1/ob ) );
    oa31_1 \U916_2_/U25/U1/Uclr  ( .x(\U916_2_/U25/U1/clr ), .a(noa), .b(a[2]), 
        .c(b[2]), .d(o[2]) );
    oaoi211_1 \U916_2_/U25/U1/Uaoi  ( .x(\U916_2_/U25/U1/ob ), .a(a[2]), .b(b
        [2]), .c(noa), .d(\U916_2_/U25/U1/clr ) );
    inv_2 \U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U916_2_/U25/U1/ob ) );
    oa31_1 \U916_3_/U25/U1/Uclr  ( .x(\U916_3_/U25/U1/clr ), .a(noa), .b(a[3]), 
        .c(b[3]), .d(o[3]) );
    oaoi211_1 \U916_3_/U25/U1/Uaoi  ( .x(\U916_3_/U25/U1/ob ), .a(a[3]), .b(b
        [3]), .c(noa), .d(\U916_3_/U25/U1/clr ) );
    inv_2 \U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U916_3_/U25/U1/ob ) );
    ao222_2 \U1148/U19/U1/U1  ( .x(o[4]), .a(noa), .b(b[4]), .c(noa), .d(o[4]), 
        .e(b[4]), .f(o[4]) );
    aoi21_1 \U1153/U11  ( .x(seta), .a(o[4]), .b(setb), .c(reset) );
    and3_3 U1 ( .x(nba), .a(bsel), .b(\noack[0] ), .c(\noack[1] ) );
endmodule


module initiator_tic ( cack, chaincommand, err, nchainresponseack, nrouteack, 
    rd, routetxreq, rrnw, a, chainresponse, col, crnw, itag, lock, nReset, 
    nchaincommandack, pred, rack, route, routetxack, seq, size, wd );
output [4:0] chaincommand;
output [1:0] err;
output [63:0] rd;
output [1:0] rrnw;
input  [63:0] a;
input  [4:0] chainresponse;
input  [5:0] col;
input  [1:0] crnw;
input  [9:0] itag;
input  [1:0] lock;
input  [1:0] pred;
input  [4:0] route;
input  [1:0] seq;
input  [3:0] size;
input  [63:0] wd;
input  nReset, nchaincommandack, rack, routetxack;
output cack, nchainresponseack, nrouteack, routetxreq;
    wire \irbh[7] , \irbh[6] , \irbh[5] , \irbh[4] , \irbh[3] , \irbh[2] , 
        \irbh[1] , \irbh[0] , \ipayload[4] , \ipayload[3] , \ipayload[2] , 
        \ipayload[1] , \ipayload[0] , \icbh[7] , \icbh[6] , \icbh[5] , 
        \icbh[4] , \icbh[3] , \icbh[2] , \icbh[1] , \icbh[0] , \cstatus[1] , 
        \cstatus[0] , \irbl[7] , \irbl[6] , \irbl[5] , \irbl[4] , \irbl[3] , 
        \irbl[2] , \irbl[1] , \irbl[0] , \rstatus[1] , \rstatus[0] , 
        \can_defer[0] , \icbl[7] , \icbl[6] , \icbl[5] , \icbl[4] , \icbl[3] , 
        \icbl[2] , \icbl[1] , \icbl[0] , nircba, nResetb, responseack, 
        rstatusack, net165, reset, tok_ack, net170, ictrlack, icmdack, 
        ncstatusack, net116, pltxreq, net115, net128, pltxack, nicba, 
        nipayloadack, \U1662/U28/U1/clr , \U1662/U28/U1/set ;
    chain_irdemuxNew_2 U1442 ( .err(err), .ncback(nircba), .rd(rd), .rnw(rrnw), 
        .status({\rstatus[1] , \rstatus[0] }), .cbh({\irbh[7] , \irbh[6] , 
        \irbh[5] , \irbh[4] , \irbh[3] , \irbh[2] , \irbh[1] , \irbh[0] }), 
        .cbl({\irbl[7] , \irbl[6] , \irbl[5] , \irbl[4] , \irbl[3] , \irbl[2] , 
        \irbl[1] , \irbl[0] }), .nReset(nResetb), .nack(responseack), 
        .statusack(rstatusack) );
    chain_fr2dr_byte_5 chain_decoder ( .nia(nchainresponseack), .oh({\irbh[7] , 
        \irbh[6] , \irbh[5] , \irbh[4] , \irbh[3] , \irbh[2] , \irbh[1] , 
        \irbh[0] }), .ol({\irbl[7] , \irbl[6] , \irbl[5] , \irbl[4] , 
        \irbl[3] , \irbl[2] , \irbl[1] , \irbl[0] }), .i(chainresponse), 
        .nReset(nResetb), .noa(nircba) );
    chain_ic_ctrl_2 cmd_ctrl ( .ack(ictrlack), .candefer(\can_defer[0] ), 
        .eop(net116), .nstatack(ncstatusack), .pltxreq(pltxreq), .routetxreq(
        routetxreq), .tok_ack(tok_ack), .accept(\cstatus[0] ), .candefer_ack({
        1'b0, \can_defer[0] }), .defer(\cstatus[1] ), .eopack(net115), .lock(
        lock), .nReset(net128), .pltxack(pltxack), .routetxack(routetxack), 
        .tok_err(err[1]), .tok_ok(err[0]) );
    chain_icmux_2 cmd_mux ( .ack(icmdack), .chainh({\icbh[7] , \icbh[6] , 
        \icbh[5] , \icbh[4] , \icbh[3] , \icbh[2] , \icbh[1] , \icbh[0] }), 
        .chainl({\icbl[7] , \icbl[6] , \icbl[5] , \icbl[4] , \icbl[3] , 
        \icbl[2] , \icbl[1] , \icbl[0] }), .sendack(pltxack), .addr(a), .col(
        col), .itag(itag), .lock(lock), .nReset(net128), .nia(nicba), .pred(
        pred), .rnw(crnw), .sendreq(pltxreq), .seq(seq), .size(size), .wd(wd)
         );
    chain_dr2fr_byte_2 U1604 ( .eop_ack(net115), .ia(nicba), .o({\ipayload[4] , 
        \ipayload[3] , \ipayload[2] , \ipayload[1] , \ipayload[0] }), .eop(
        net116), .ih({\icbh[7] , \icbh[6] , \icbh[5] , \icbh[4] , \icbh[3] , 
        \icbh[2] , \icbh[1] , \icbh[0] }), .il({\icbl[7] , \icbl[6] , 
        \icbl[5] , \icbl[4] , \icbl[3] , \icbl[2] , \icbl[1] , \icbl[0] }), 
        .nReset(net128), .noa(nipayloadack) );
    chain_mergepackets_2 U1605 ( .naa(nrouteack), .nba(nipayloadack), .o(
        chaincommand), .a(route), .b({\ipayload[4] , \ipayload[3] , 
        \ipayload[2] , \ipayload[1] , \ipayload[0] }), .nReset(net128), .noa(
        nchaincommandack) );
    and2_1 U1676 ( .x(cack), .a(net170), .b(nResetb) );
    inv_4 \U1643/U3  ( .x(net128), .a(reset) );
    or2_4 \U1660/U12  ( .x(net165), .a(\cstatus[0] ), .b(\cstatus[1] ) );
    or2_1 \U1661/U12  ( .x(rstatusack), .a(net165), .b(reset) );
    ao222_2 \status_pipe_0_/U19/U1/U1  ( .x(\cstatus[0] ), .a(\rstatus[0] ), 
        .b(ncstatusack), .c(\rstatus[0] ), .d(\cstatus[0] ), .e(ncstatusack), 
        .f(\cstatus[0] ) );
    ao222_2 \status_pipe_1_/U19/U1/U1  ( .x(\cstatus[1] ), .a(\rstatus[1] ), 
        .b(ncstatusack), .c(\rstatus[1] ), .d(\cstatus[1] ), .e(ncstatusack), 
        .f(\cstatus[1] ) );
    ao222_1 \U1609/U18/U1/U1  ( .x(net170), .a(ictrlack), .b(icmdack), .c(
        ictrlack), .d(net170), .e(icmdack), .f(net170) );
    aoai211_1 \U1662/U28/U1/U1  ( .x(\U1662/U28/U1/clr ), .a(rack), .b(nResetb
        ), .c(tok_ack), .d(responseack) );
    nand3_1 \U1662/U28/U1/U2  ( .x(\U1662/U28/U1/set ), .a(tok_ack), .b(rack), 
        .c(nResetb) );
    nand2_2 \U1662/U28/U1/U3  ( .x(responseack), .a(\U1662/U28/U1/clr ), .b(
        \U1662/U28/U1/set ) );
    inv_2 U1 ( .x(reset), .a(nResetb) );
    buf_3 U2 ( .x(nResetb), .a(nReset) );
endmodule


module matched_delay_m2cp_com_tic ( x, a );
input  a;
output x;
    wire n2;
    buf_1 I1 ( .x(n2), .a(a) );
    buf_16 U1 ( .x(x), .a(n2) );
endmodule


module matched_delay_m2cp_resp_tic ( x, a );
input  a;
output x;
    assign x = a;
endmodule


module sr2dr_word_4 ( i, req, h, l );
input  [31:0] i;
output [31:0] h;
output [31:0] l;
input  req;
    wire \U31/nl , \U31/ni , \U31/nh , \U30/nl , \U30/ni , \U30/nh , \U29/nl , 
        \U29/ni , \U29/nh , \U28/nl , \U28/ni , \U28/nh , \U27/nl , \U27/ni , 
        \U27/nh , \U26/nl , \U26/ni , \U26/nh , \U25/nl , \U25/ni , \U25/nh , 
        \U24/nl , \U24/ni , \U24/nh , \U23/nl , \U23/ni , \U23/nh , \U22/nl , 
        \U22/ni , \U22/nh , \U21/nl , \U21/ni , \U21/nh , \U20/nl , \U20/ni , 
        \U20/nh , \U19/nl , \U19/ni , \U19/nh , \U18/nl , \U18/ni , \U18/nh , 
        \U17/nl , \U17/ni , \U17/nh , \U16/nl , \U16/ni , \U16/nh , \U15/nl , 
        \U15/ni , \U15/nh , \U14/nl , \U14/ni , \U14/nh , \U13/nl , \U13/ni , 
        \U13/nh , \U12/nl , \U12/ni , \U12/nh , \U11/nl , \U11/ni , \U11/nh , 
        \U10/nl , \U10/ni , \U10/nh , \U9/nl , \U9/ni , \U9/nh , \U8/nl , 
        \U8/ni , \U8/nh , \U7/nl , \U7/ni , \U7/nh , \U6/nl , \U6/ni , \U6/nh , 
        \U5/nl , \U5/ni , \U5/nh , \U4/nl , \U4/ni , \U4/nh , \U3/nl , \U3/ni , 
        \U3/nh , \U2/nl , \U2/ni , \U2/nh , \U1/nl , \U1/ni , \U1/nh , \U0/nl , 
        \U0/ni , \U0/nh , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
    inv_1 \U31/Uii  ( .x(\U31/ni ), .a(i[31]) );
    inv_1 \U31/Uih  ( .x(\U31/nh ), .a(h[31]) );
    inv_1 \U31/Uil  ( .x(\U31/nl ), .a(l[31]) );
    ao23_1 \U31/Ucl/U1/U1  ( .x(l[31]), .a(n9), .b(l[31]), .c(n1), .d(\U31/ni 
        ), .e(\U31/nh ) );
    ao23_1 \U31/Uch/U1/U1  ( .x(h[31]), .a(n9), .b(h[31]), .c(n2), .d(i[31]), 
        .e(\U31/nl ) );
    inv_1 \U30/Uii  ( .x(\U30/ni ), .a(i[30]) );
    inv_1 \U30/Uih  ( .x(\U30/nh ), .a(h[30]) );
    inv_1 \U30/Uil  ( .x(\U30/nl ), .a(l[30]) );
    ao23_1 \U30/Ucl/U1/U1  ( .x(l[30]), .a(n8), .b(l[30]), .c(n1), .d(\U30/ni 
        ), .e(\U30/nh ) );
    ao23_1 \U30/Uch/U1/U1  ( .x(h[30]), .a(n8), .b(h[30]), .c(n1), .d(i[30]), 
        .e(\U30/nl ) );
    inv_1 \U29/Uii  ( .x(\U29/ni ), .a(i[29]) );
    inv_1 \U29/Uih  ( .x(\U29/nh ), .a(h[29]) );
    inv_1 \U29/Uil  ( .x(\U29/nl ), .a(l[29]) );
    ao23_1 \U29/Ucl/U1/U1  ( .x(l[29]), .a(n8), .b(l[29]), .c(n1), .d(\U29/ni 
        ), .e(\U29/nh ) );
    ao23_1 \U29/Uch/U1/U1  ( .x(h[29]), .a(n8), .b(h[29]), .c(n2), .d(i[29]), 
        .e(\U29/nl ) );
    inv_1 \U28/Uii  ( .x(\U28/ni ), .a(i[28]) );
    inv_1 \U28/Uih  ( .x(\U28/nh ), .a(h[28]) );
    inv_1 \U28/Uil  ( .x(\U28/nl ), .a(l[28]) );
    ao23_1 \U28/Ucl/U1/U1  ( .x(l[28]), .a(n8), .b(l[28]), .c(n2), .d(\U28/ni 
        ), .e(\U28/nh ) );
    ao23_1 \U28/Uch/U1/U1  ( .x(h[28]), .a(n8), .b(h[28]), .c(n2), .d(i[28]), 
        .e(\U28/nl ) );
    inv_1 \U27/Uii  ( .x(\U27/ni ), .a(i[27]) );
    inv_1 \U27/Uih  ( .x(\U27/nh ), .a(h[27]) );
    inv_1 \U27/Uil  ( .x(\U27/nl ), .a(l[27]) );
    ao23_1 \U27/Ucl/U1/U1  ( .x(l[27]), .a(n8), .b(l[27]), .c(n2), .d(\U27/ni 
        ), .e(\U27/nh ) );
    ao23_1 \U27/Uch/U1/U1  ( .x(h[27]), .a(n8), .b(h[27]), .c(n2), .d(i[27]), 
        .e(\U27/nl ) );
    inv_1 \U26/Uii  ( .x(\U26/ni ), .a(i[26]) );
    inv_1 \U26/Uih  ( .x(\U26/nh ), .a(h[26]) );
    inv_1 \U26/Uil  ( .x(\U26/nl ), .a(l[26]) );
    ao23_1 \U26/Ucl/U1/U1  ( .x(l[26]), .a(n7), .b(l[26]), .c(n2), .d(\U26/ni 
        ), .e(\U26/nh ) );
    ao23_1 \U26/Uch/U1/U1  ( .x(h[26]), .a(n7), .b(h[26]), .c(n4), .d(i[26]), 
        .e(\U26/nl ) );
    inv_1 \U25/Uii  ( .x(\U25/ni ), .a(i[25]) );
    inv_1 \U25/Uih  ( .x(\U25/nh ), .a(h[25]) );
    inv_1 \U25/Uil  ( .x(\U25/nl ), .a(l[25]) );
    ao23_1 \U25/Ucl/U1/U1  ( .x(l[25]), .a(n7), .b(l[25]), .c(n4), .d(\U25/ni 
        ), .e(\U25/nh ) );
    ao23_1 \U25/Uch/U1/U1  ( .x(h[25]), .a(n7), .b(h[25]), .c(n4), .d(i[25]), 
        .e(\U25/nl ) );
    inv_1 \U24/Uii  ( .x(\U24/ni ), .a(i[24]) );
    inv_1 \U24/Uih  ( .x(\U24/nh ), .a(h[24]) );
    inv_1 \U24/Uil  ( .x(\U24/nl ), .a(l[24]) );
    ao23_1 \U24/Ucl/U1/U1  ( .x(l[24]), .a(n7), .b(l[24]), .c(n4), .d(\U24/ni 
        ), .e(\U24/nh ) );
    ao23_1 \U24/Uch/U1/U1  ( .x(h[24]), .a(n7), .b(h[24]), .c(n4), .d(i[24]), 
        .e(\U24/nl ) );
    inv_1 \U23/Uii  ( .x(\U23/ni ), .a(i[23]) );
    inv_1 \U23/Uih  ( .x(\U23/nh ), .a(h[23]) );
    inv_1 \U23/Uil  ( .x(\U23/nl ), .a(l[23]) );
    ao23_1 \U23/Ucl/U1/U1  ( .x(l[23]), .a(n7), .b(l[23]), .c(n3), .d(\U23/ni 
        ), .e(\U23/nh ) );
    ao23_1 \U23/Uch/U1/U1  ( .x(h[23]), .a(n7), .b(h[23]), .c(n3), .d(i[23]), 
        .e(\U23/nl ) );
    inv_1 \U22/Uii  ( .x(\U22/ni ), .a(i[22]) );
    inv_1 \U22/Uih  ( .x(\U22/nh ), .a(h[22]) );
    inv_1 \U22/Uil  ( .x(\U22/nl ), .a(l[22]) );
    ao23_1 \U22/Ucl/U1/U1  ( .x(l[22]), .a(n6), .b(l[22]), .c(n3), .d(\U22/ni 
        ), .e(\U22/nh ) );
    ao23_1 \U22/Uch/U1/U1  ( .x(h[22]), .a(n6), .b(h[22]), .c(n3), .d(i[22]), 
        .e(\U22/nl ) );
    inv_1 \U21/Uii  ( .x(\U21/ni ), .a(i[21]) );
    inv_1 \U21/Uih  ( .x(\U21/nh ), .a(h[21]) );
    inv_1 \U21/Uil  ( .x(\U21/nl ), .a(l[21]) );
    ao23_1 \U21/Ucl/U1/U1  ( .x(l[21]), .a(n6), .b(l[21]), .c(n3), .d(\U21/ni 
        ), .e(\U21/nh ) );
    ao23_1 \U21/Uch/U1/U1  ( .x(h[21]), .a(n6), .b(h[21]), .c(n3), .d(i[21]), 
        .e(\U21/nl ) );
    inv_1 \U20/Uii  ( .x(\U20/ni ), .a(i[20]) );
    inv_1 \U20/Uih  ( .x(\U20/nh ), .a(h[20]) );
    inv_1 \U20/Uil  ( .x(\U20/nl ), .a(l[20]) );
    ao23_1 \U20/Ucl/U1/U1  ( .x(l[20]), .a(n6), .b(l[20]), .c(n5), .d(\U20/ni 
        ), .e(\U20/nh ) );
    ao23_1 \U20/Uch/U1/U1  ( .x(h[20]), .a(n6), .b(h[20]), .c(n4), .d(i[20]), 
        .e(\U20/nl ) );
    inv_1 \U19/Uii  ( .x(\U19/ni ), .a(i[19]) );
    inv_1 \U19/Uih  ( .x(\U19/nh ), .a(h[19]) );
    inv_1 \U19/Uil  ( .x(\U19/nl ), .a(l[19]) );
    ao23_1 \U19/Ucl/U1/U1  ( .x(l[19]), .a(n6), .b(l[19]), .c(n4), .d(\U19/ni 
        ), .e(\U19/nh ) );
    ao23_1 \U19/Uch/U1/U1  ( .x(h[19]), .a(n6), .b(h[19]), .c(n4), .d(i[19]), 
        .e(\U19/nl ) );
    inv_1 \U18/Uii  ( .x(\U18/ni ), .a(i[18]) );
    inv_1 \U18/Uih  ( .x(\U18/nh ), .a(h[18]) );
    inv_1 \U18/Uil  ( .x(\U18/nl ), .a(l[18]) );
    ao23_1 \U18/Ucl/U1/U1  ( .x(l[18]), .a(n5), .b(l[18]), .c(n5), .d(\U18/ni 
        ), .e(\U18/nh ) );
    ao23_1 \U18/Uch/U1/U1  ( .x(h[18]), .a(n5), .b(h[18]), .c(n5), .d(i[18]), 
        .e(\U18/nl ) );
    inv_1 \U17/Uii  ( .x(\U17/ni ), .a(i[17]) );
    inv_1 \U17/Uih  ( .x(\U17/nh ), .a(h[17]) );
    inv_1 \U17/Uil  ( .x(\U17/nl ), .a(l[17]) );
    ao23_1 \U17/Ucl/U1/U1  ( .x(l[17]), .a(n6), .b(l[17]), .c(n5), .d(\U17/ni 
        ), .e(\U17/nh ) );
    ao23_1 \U17/Uch/U1/U1  ( .x(h[17]), .a(n7), .b(h[17]), .c(n4), .d(i[17]), 
        .e(\U17/nl ) );
    inv_1 \U16/Uii  ( .x(\U16/ni ), .a(i[16]) );
    inv_1 \U16/Uih  ( .x(\U16/nh ), .a(h[16]) );
    inv_1 \U16/Uil  ( .x(\U16/nl ), .a(l[16]) );
    ao23_1 \U16/Ucl/U1/U1  ( .x(l[16]), .a(n9), .b(l[16]), .c(n3), .d(\U16/ni 
        ), .e(\U16/nh ) );
    ao23_1 \U16/Uch/U1/U1  ( .x(h[16]), .a(n9), .b(h[16]), .c(n1), .d(i[16]), 
        .e(\U16/nl ) );
    inv_1 \U15/Uii  ( .x(\U15/ni ), .a(i[15]) );
    inv_1 \U15/Uih  ( .x(\U15/nh ), .a(h[15]) );
    inv_1 \U15/Uil  ( .x(\U15/nl ), .a(l[15]) );
    ao23_1 \U15/Ucl/U1/U1  ( .x(l[15]), .a(n8), .b(l[15]), .c(n1), .d(\U15/ni 
        ), .e(\U15/nh ) );
    ao23_1 \U15/Uch/U1/U1  ( .x(h[15]), .a(n7), .b(h[15]), .c(n1), .d(i[15]), 
        .e(\U15/nl ) );
    inv_1 \U14/Uii  ( .x(\U14/ni ), .a(i[14]) );
    inv_1 \U14/Uih  ( .x(\U14/nh ), .a(h[14]) );
    inv_1 \U14/Uil  ( .x(\U14/nl ), .a(l[14]) );
    ao23_1 \U14/Ucl/U1/U1  ( .x(l[14]), .a(n6), .b(l[14]), .c(n1), .d(\U14/ni 
        ), .e(\U14/nh ) );
    ao23_1 \U14/Uch/U1/U1  ( .x(h[14]), .a(n6), .b(h[14]), .c(n3), .d(i[14]), 
        .e(\U14/nl ) );
    inv_1 \U13/Uii  ( .x(\U13/ni ), .a(i[13]) );
    inv_1 \U13/Uih  ( .x(\U13/nh ), .a(h[13]) );
    inv_1 \U13/Uil  ( .x(\U13/nl ), .a(l[13]) );
    ao23_1 \U13/Ucl/U1/U1  ( .x(l[13]), .a(n6), .b(l[13]), .c(n4), .d(\U13/ni 
        ), .e(\U13/nh ) );
    ao23_1 \U13/Uch/U1/U1  ( .x(h[13]), .a(n6), .b(h[13]), .c(n4), .d(i[13]), 
        .e(\U13/nl ) );
    inv_1 \U12/Uii  ( .x(\U12/ni ), .a(i[12]) );
    inv_1 \U12/Uih  ( .x(\U12/nh ), .a(h[12]) );
    inv_1 \U12/Uil  ( .x(\U12/nl ), .a(l[12]) );
    ao23_1 \U12/Ucl/U1/U1  ( .x(l[12]), .a(n5), .b(l[12]), .c(n4), .d(\U12/ni 
        ), .e(\U12/nh ) );
    ao23_1 \U12/Uch/U1/U1  ( .x(h[12]), .a(n5), .b(h[12]), .c(n4), .d(i[12]), 
        .e(\U12/nl ) );
    inv_1 \U11/Uii  ( .x(\U11/ni ), .a(i[11]) );
    inv_1 \U11/Uih  ( .x(\U11/nh ), .a(h[11]) );
    inv_1 \U11/Uil  ( .x(\U11/nl ), .a(l[11]) );
    ao23_1 \U11/Ucl/U1/U1  ( .x(l[11]), .a(n5), .b(l[11]), .c(n4), .d(\U11/ni 
        ), .e(\U11/nh ) );
    ao23_1 \U11/Uch/U1/U1  ( .x(h[11]), .a(n5), .b(h[11]), .c(n4), .d(i[11]), 
        .e(\U11/nl ) );
    inv_1 \U10/Uii  ( .x(\U10/ni ), .a(i[10]) );
    inv_1 \U10/Uih  ( .x(\U10/nh ), .a(h[10]) );
    inv_1 \U10/Uil  ( .x(\U10/nl ), .a(l[10]) );
    ao23_1 \U10/Ucl/U1/U1  ( .x(l[10]), .a(n5), .b(l[10]), .c(n3), .d(\U10/ni 
        ), .e(\U10/nh ) );
    ao23_1 \U10/Uch/U1/U1  ( .x(h[10]), .a(n5), .b(h[10]), .c(n3), .d(i[10]), 
        .e(\U10/nl ) );
    inv_1 \U9/Uii  ( .x(\U9/ni ), .a(i[9]) );
    inv_1 \U9/Uih  ( .x(\U9/nh ), .a(h[9]) );
    inv_1 \U9/Uil  ( .x(\U9/nl ), .a(l[9]) );
    ao23_1 \U9/Ucl/U1/U1  ( .x(l[9]), .a(n5), .b(l[9]), .c(n3), .d(\U9/ni ), 
        .e(\U9/nh ) );
    ao23_1 \U9/Uch/U1/U1  ( .x(h[9]), .a(n5), .b(h[9]), .c(n3), .d(i[9]), .e(
        \U9/nl ) );
    inv_1 \U8/Uii  ( .x(\U8/ni ), .a(i[8]) );
    inv_1 \U8/Uih  ( .x(\U8/nh ), .a(h[8]) );
    inv_1 \U8/Uil  ( .x(\U8/nl ), .a(l[8]) );
    ao23_1 \U8/Ucl/U1/U1  ( .x(l[8]), .a(n5), .b(l[8]), .c(n3), .d(\U8/ni ), 
        .e(\U8/nh ) );
    ao23_1 \U8/Uch/U1/U1  ( .x(h[8]), .a(n5), .b(h[8]), .c(n3), .d(i[8]), .e(
        \U8/nl ) );
    inv_1 \U7/Uii  ( .x(\U7/ni ), .a(i[7]) );
    inv_1 \U7/Uih  ( .x(\U7/nh ), .a(h[7]) );
    inv_1 \U7/Uil  ( .x(\U7/nl ), .a(l[7]) );
    ao23_1 \U7/Ucl/U1/U1  ( .x(l[7]), .a(n7), .b(l[7]), .c(n3), .d(\U7/ni ), 
        .e(\U7/nh ) );
    ao23_1 \U7/Uch/U1/U1  ( .x(h[7]), .a(n7), .b(h[7]), .c(n2), .d(i[7]), .e(
        \U7/nl ) );
    inv_1 \U6/Uii  ( .x(\U6/ni ), .a(i[6]) );
    inv_1 \U6/Uih  ( .x(\U6/nh ), .a(h[6]) );
    inv_1 \U6/Uil  ( .x(\U6/nl ), .a(l[6]) );
    ao23_1 \U6/Ucl/U1/U1  ( .x(l[6]), .a(n7), .b(l[6]), .c(n2), .d(\U6/ni ), 
        .e(\U6/nh ) );
    ao23_1 \U6/Uch/U1/U1  ( .x(h[6]), .a(n7), .b(h[6]), .c(n2), .d(i[6]), .e(
        \U6/nl ) );
    inv_1 \U5/Uii  ( .x(\U5/ni ), .a(i[5]) );
    inv_1 \U5/Uih  ( .x(\U5/nh ), .a(h[5]) );
    inv_1 \U5/Uil  ( .x(\U5/nl ), .a(l[5]) );
    ao23_1 \U5/Ucl/U1/U1  ( .x(l[5]), .a(n7), .b(l[5]), .c(n2), .d(\U5/ni ), 
        .e(\U5/nh ) );
    ao23_1 \U5/Uch/U1/U1  ( .x(h[5]), .a(n7), .b(h[5]), .c(n2), .d(i[5]), .e(
        \U5/nl ) );
    inv_1 \U4/Uii  ( .x(\U4/ni ), .a(i[4]) );
    inv_1 \U4/Uih  ( .x(\U4/nh ), .a(h[4]) );
    inv_1 \U4/Uil  ( .x(\U4/nl ), .a(l[4]) );
    ao23_1 \U4/Ucl/U1/U1  ( .x(l[4]), .a(n6), .b(l[4]), .c(n2), .d(\U4/ni ), 
        .e(\U4/nh ) );
    ao23_1 \U4/Uch/U1/U1  ( .x(h[4]), .a(n6), .b(h[4]), .c(n2), .d(i[4]), .e(
        \U4/nl ) );
    inv_1 \U3/Uii  ( .x(\U3/ni ), .a(i[3]) );
    inv_1 \U3/Uih  ( .x(\U3/nh ), .a(h[3]) );
    inv_1 \U3/Uil  ( .x(\U3/nl ), .a(l[3]) );
    ao23_1 \U3/Ucl/U1/U1  ( .x(l[3]), .a(n6), .b(l[3]), .c(n2), .d(\U3/ni ), 
        .e(\U3/nh ) );
    ao23_1 \U3/Uch/U1/U1  ( .x(h[3]), .a(n8), .b(h[3]), .c(n1), .d(i[3]), .e(
        \U3/nl ) );
    inv_1 \U2/Uii  ( .x(\U2/ni ), .a(i[2]) );
    inv_1 \U2/Uih  ( .x(\U2/nh ), .a(h[2]) );
    inv_1 \U2/Uil  ( .x(\U2/nl ), .a(l[2]) );
    ao23_1 \U2/Ucl/U1/U1  ( .x(l[2]), .a(n8), .b(l[2]), .c(n1), .d(\U2/ni ), 
        .e(\U2/nh ) );
    ao23_1 \U2/Uch/U1/U1  ( .x(h[2]), .a(n8), .b(h[2]), .c(n1), .d(i[2]), .e(
        \U2/nl ) );
    inv_1 \U1/Uii  ( .x(\U1/ni ), .a(i[1]) );
    inv_1 \U1/Uih  ( .x(\U1/nh ), .a(h[1]) );
    inv_1 \U1/Uil  ( .x(\U1/nl ), .a(l[1]) );
    ao23_1 \U1/Ucl/U1/U1  ( .x(l[1]), .a(n8), .b(l[1]), .c(n1), .d(\U1/ni ), 
        .e(\U1/nh ) );
    ao23_1 \U1/Uch/U1/U1  ( .x(h[1]), .a(n8), .b(h[1]), .c(n1), .d(i[1]), .e(
        \U1/nl ) );
    inv_1 \U0/Uii  ( .x(\U0/ni ), .a(i[0]) );
    inv_1 \U0/Uih  ( .x(\U0/nh ), .a(h[0]) );
    inv_1 \U0/Uil  ( .x(\U0/nl ), .a(l[0]) );
    ao23_1 \U0/Ucl/U1/U1  ( .x(l[0]), .a(n8), .b(l[0]), .c(n1), .d(\U0/ni ), 
        .e(\U0/nh ) );
    ao23_1 \U0/Uch/U1/U1  ( .x(h[0]), .a(n8), .b(h[0]), .c(n1), .d(i[0]), .e(
        \U0/nl ) );
    buf_16 U1 ( .x(n1), .a(n12) );
    buf_16 U2 ( .x(n2), .a(n12) );
    buf_16 U3 ( .x(n3), .a(n12) );
    buf_16 U4 ( .x(n4), .a(n11) );
    buf_16 U5 ( .x(n5), .a(n11) );
    buf_16 U6 ( .x(n6), .a(n11) );
    buf_16 U7 ( .x(n7), .a(n10) );
    buf_16 U8 ( .x(n8), .a(n10) );
    buf_16 U9 ( .x(n9), .a(n10) );
    buf_16 U10 ( .x(n10), .a(req) );
    buf_16 U11 ( .x(n11), .a(req) );
    buf_16 U12 ( .x(n12), .a(req) );
endmodule


module sr2dr_word_5 ( i, req, h, l );
input  [31:0] i;
output [31:0] h;
output [31:0] l;
input  req;
    wire \U31/nl , \U31/ni , \U31/nh , \U30/nl , \U30/ni , \U30/nh , \U29/nl , 
        \U29/ni , \U29/nh , \U28/nl , \U28/ni , \U28/nh , \U27/nl , \U27/ni , 
        \U27/nh , \U26/nl , \U26/ni , \U26/nh , \U25/nl , \U25/ni , \U25/nh , 
        \U24/nl , \U24/ni , \U24/nh , \U23/nl , \U23/ni , \U23/nh , \U22/nl , 
        \U22/ni , \U22/nh , \U21/nl , \U21/ni , \U21/nh , \U20/nl , \U20/ni , 
        \U20/nh , \U19/nl , \U19/ni , \U19/nh , \U18/nl , \U18/ni , \U18/nh , 
        \U17/nl , \U17/ni , \U17/nh , \U16/nl , \U16/ni , \U16/nh , \U15/nl , 
        \U15/ni , \U15/nh , \U14/nl , \U14/ni , \U14/nh , \U13/nl , \U13/ni , 
        \U13/nh , \U12/nl , \U12/ni , \U12/nh , \U11/nl , \U11/ni , \U11/nh , 
        \U10/nl , \U10/ni , \U10/nh , \U9/nl , \U9/ni , \U9/nh , \U8/nl , 
        \U8/ni , \U8/nh , \U7/nl , \U7/ni , \U7/nh , \U6/nl , \U6/ni , \U6/nh , 
        \U5/nl , \U5/ni , \U5/nh , \U4/nl , \U4/ni , \U4/nh , \U3/nl , \U3/ni , 
        \U3/nh , \U2/nl , \U2/ni , \U2/nh , \U1/nl , \U1/ni , \U1/nh , \U0/nl , 
        \U0/ni , \U0/nh , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
    inv_1 \U31/Uii  ( .x(\U31/ni ), .a(i[31]) );
    inv_1 \U31/Uih  ( .x(\U31/nh ), .a(h[31]) );
    inv_1 \U31/Uil  ( .x(\U31/nl ), .a(l[31]) );
    ao23_1 \U31/Ucl/U1/U1  ( .x(l[31]), .a(n9), .b(l[31]), .c(n1), .d(\U31/ni 
        ), .e(\U31/nh ) );
    ao23_1 \U31/Uch/U1/U1  ( .x(h[31]), .a(n9), .b(h[31]), .c(n2), .d(i[31]), 
        .e(\U31/nl ) );
    inv_1 \U30/Uii  ( .x(\U30/ni ), .a(i[30]) );
    inv_1 \U30/Uih  ( .x(\U30/nh ), .a(h[30]) );
    inv_1 \U30/Uil  ( .x(\U30/nl ), .a(l[30]) );
    ao23_1 \U30/Ucl/U1/U1  ( .x(l[30]), .a(n8), .b(l[30]), .c(n1), .d(\U30/ni 
        ), .e(\U30/nh ) );
    ao23_1 \U30/Uch/U1/U1  ( .x(h[30]), .a(n8), .b(h[30]), .c(n1), .d(i[30]), 
        .e(\U30/nl ) );
    inv_1 \U29/Uii  ( .x(\U29/ni ), .a(i[29]) );
    inv_1 \U29/Uih  ( .x(\U29/nh ), .a(h[29]) );
    inv_1 \U29/Uil  ( .x(\U29/nl ), .a(l[29]) );
    ao23_1 \U29/Ucl/U1/U1  ( .x(l[29]), .a(n8), .b(l[29]), .c(n1), .d(\U29/ni 
        ), .e(\U29/nh ) );
    ao23_1 \U29/Uch/U1/U1  ( .x(h[29]), .a(n8), .b(h[29]), .c(n2), .d(i[29]), 
        .e(\U29/nl ) );
    inv_1 \U28/Uii  ( .x(\U28/ni ), .a(i[28]) );
    inv_1 \U28/Uih  ( .x(\U28/nh ), .a(h[28]) );
    inv_1 \U28/Uil  ( .x(\U28/nl ), .a(l[28]) );
    ao23_1 \U28/Ucl/U1/U1  ( .x(l[28]), .a(n8), .b(l[28]), .c(n2), .d(\U28/ni 
        ), .e(\U28/nh ) );
    ao23_1 \U28/Uch/U1/U1  ( .x(h[28]), .a(n8), .b(h[28]), .c(n2), .d(i[28]), 
        .e(\U28/nl ) );
    inv_1 \U27/Uii  ( .x(\U27/ni ), .a(i[27]) );
    inv_1 \U27/Uih  ( .x(\U27/nh ), .a(h[27]) );
    inv_1 \U27/Uil  ( .x(\U27/nl ), .a(l[27]) );
    ao23_1 \U27/Ucl/U1/U1  ( .x(l[27]), .a(n8), .b(l[27]), .c(n2), .d(\U27/ni 
        ), .e(\U27/nh ) );
    ao23_1 \U27/Uch/U1/U1  ( .x(h[27]), .a(n8), .b(h[27]), .c(n2), .d(i[27]), 
        .e(\U27/nl ) );
    inv_1 \U26/Uii  ( .x(\U26/ni ), .a(i[26]) );
    inv_1 \U26/Uih  ( .x(\U26/nh ), .a(h[26]) );
    inv_1 \U26/Uil  ( .x(\U26/nl ), .a(l[26]) );
    ao23_1 \U26/Ucl/U1/U1  ( .x(l[26]), .a(n7), .b(l[26]), .c(n2), .d(\U26/ni 
        ), .e(\U26/nh ) );
    ao23_1 \U26/Uch/U1/U1  ( .x(h[26]), .a(n7), .b(h[26]), .c(n4), .d(i[26]), 
        .e(\U26/nl ) );
    inv_1 \U25/Uii  ( .x(\U25/ni ), .a(i[25]) );
    inv_1 \U25/Uih  ( .x(\U25/nh ), .a(h[25]) );
    inv_1 \U25/Uil  ( .x(\U25/nl ), .a(l[25]) );
    ao23_1 \U25/Ucl/U1/U1  ( .x(l[25]), .a(n7), .b(l[25]), .c(n4), .d(\U25/ni 
        ), .e(\U25/nh ) );
    ao23_1 \U25/Uch/U1/U1  ( .x(h[25]), .a(n7), .b(h[25]), .c(n4), .d(i[25]), 
        .e(\U25/nl ) );
    inv_1 \U24/Uii  ( .x(\U24/ni ), .a(i[24]) );
    inv_1 \U24/Uih  ( .x(\U24/nh ), .a(h[24]) );
    inv_1 \U24/Uil  ( .x(\U24/nl ), .a(l[24]) );
    ao23_1 \U24/Ucl/U1/U1  ( .x(l[24]), .a(n7), .b(l[24]), .c(n4), .d(\U24/ni 
        ), .e(\U24/nh ) );
    ao23_1 \U24/Uch/U1/U1  ( .x(h[24]), .a(n7), .b(h[24]), .c(n4), .d(i[24]), 
        .e(\U24/nl ) );
    inv_1 \U23/Uii  ( .x(\U23/ni ), .a(i[23]) );
    inv_1 \U23/Uih  ( .x(\U23/nh ), .a(h[23]) );
    inv_1 \U23/Uil  ( .x(\U23/nl ), .a(l[23]) );
    ao23_1 \U23/Ucl/U1/U1  ( .x(l[23]), .a(n7), .b(l[23]), .c(n3), .d(\U23/ni 
        ), .e(\U23/nh ) );
    ao23_1 \U23/Uch/U1/U1  ( .x(h[23]), .a(n7), .b(h[23]), .c(n3), .d(i[23]), 
        .e(\U23/nl ) );
    inv_1 \U22/Uii  ( .x(\U22/ni ), .a(i[22]) );
    inv_1 \U22/Uih  ( .x(\U22/nh ), .a(h[22]) );
    inv_1 \U22/Uil  ( .x(\U22/nl ), .a(l[22]) );
    ao23_1 \U22/Ucl/U1/U1  ( .x(l[22]), .a(n6), .b(l[22]), .c(n3), .d(\U22/ni 
        ), .e(\U22/nh ) );
    ao23_1 \U22/Uch/U1/U1  ( .x(h[22]), .a(n6), .b(h[22]), .c(n3), .d(i[22]), 
        .e(\U22/nl ) );
    inv_1 \U21/Uii  ( .x(\U21/ni ), .a(i[21]) );
    inv_1 \U21/Uih  ( .x(\U21/nh ), .a(h[21]) );
    inv_1 \U21/Uil  ( .x(\U21/nl ), .a(l[21]) );
    ao23_1 \U21/Ucl/U1/U1  ( .x(l[21]), .a(n6), .b(l[21]), .c(n3), .d(\U21/ni 
        ), .e(\U21/nh ) );
    ao23_1 \U21/Uch/U1/U1  ( .x(h[21]), .a(n6), .b(h[21]), .c(n3), .d(i[21]), 
        .e(\U21/nl ) );
    inv_1 \U20/Uii  ( .x(\U20/ni ), .a(i[20]) );
    inv_1 \U20/Uih  ( .x(\U20/nh ), .a(h[20]) );
    inv_1 \U20/Uil  ( .x(\U20/nl ), .a(l[20]) );
    ao23_1 \U20/Ucl/U1/U1  ( .x(l[20]), .a(n6), .b(l[20]), .c(n5), .d(\U20/ni 
        ), .e(\U20/nh ) );
    ao23_1 \U20/Uch/U1/U1  ( .x(h[20]), .a(n6), .b(h[20]), .c(n4), .d(i[20]), 
        .e(\U20/nl ) );
    inv_1 \U19/Uii  ( .x(\U19/ni ), .a(i[19]) );
    inv_1 \U19/Uih  ( .x(\U19/nh ), .a(h[19]) );
    inv_1 \U19/Uil  ( .x(\U19/nl ), .a(l[19]) );
    ao23_1 \U19/Ucl/U1/U1  ( .x(l[19]), .a(n6), .b(l[19]), .c(n4), .d(\U19/ni 
        ), .e(\U19/nh ) );
    ao23_1 \U19/Uch/U1/U1  ( .x(h[19]), .a(n6), .b(h[19]), .c(n4), .d(i[19]), 
        .e(\U19/nl ) );
    inv_1 \U18/Uii  ( .x(\U18/ni ), .a(i[18]) );
    inv_1 \U18/Uih  ( .x(\U18/nh ), .a(h[18]) );
    inv_1 \U18/Uil  ( .x(\U18/nl ), .a(l[18]) );
    ao23_1 \U18/Ucl/U1/U1  ( .x(l[18]), .a(n5), .b(l[18]), .c(n5), .d(\U18/ni 
        ), .e(\U18/nh ) );
    ao23_1 \U18/Uch/U1/U1  ( .x(h[18]), .a(n5), .b(h[18]), .c(n5), .d(i[18]), 
        .e(\U18/nl ) );
    inv_1 \U17/Uii  ( .x(\U17/ni ), .a(i[17]) );
    inv_1 \U17/Uih  ( .x(\U17/nh ), .a(h[17]) );
    inv_1 \U17/Uil  ( .x(\U17/nl ), .a(l[17]) );
    ao23_1 \U17/Ucl/U1/U1  ( .x(l[17]), .a(n6), .b(l[17]), .c(n5), .d(\U17/ni 
        ), .e(\U17/nh ) );
    ao23_1 \U17/Uch/U1/U1  ( .x(h[17]), .a(n7), .b(h[17]), .c(n4), .d(i[17]), 
        .e(\U17/nl ) );
    inv_1 \U16/Uii  ( .x(\U16/ni ), .a(i[16]) );
    inv_1 \U16/Uih  ( .x(\U16/nh ), .a(h[16]) );
    inv_1 \U16/Uil  ( .x(\U16/nl ), .a(l[16]) );
    ao23_1 \U16/Ucl/U1/U1  ( .x(l[16]), .a(n9), .b(l[16]), .c(n3), .d(\U16/ni 
        ), .e(\U16/nh ) );
    ao23_1 \U16/Uch/U1/U1  ( .x(h[16]), .a(n9), .b(h[16]), .c(n1), .d(i[16]), 
        .e(\U16/nl ) );
    inv_1 \U15/Uii  ( .x(\U15/ni ), .a(i[15]) );
    inv_1 \U15/Uih  ( .x(\U15/nh ), .a(h[15]) );
    inv_1 \U15/Uil  ( .x(\U15/nl ), .a(l[15]) );
    ao23_1 \U15/Ucl/U1/U1  ( .x(l[15]), .a(n8), .b(l[15]), .c(n1), .d(\U15/ni 
        ), .e(\U15/nh ) );
    ao23_1 \U15/Uch/U1/U1  ( .x(h[15]), .a(n7), .b(h[15]), .c(n1), .d(i[15]), 
        .e(\U15/nl ) );
    inv_1 \U14/Uii  ( .x(\U14/ni ), .a(i[14]) );
    inv_1 \U14/Uih  ( .x(\U14/nh ), .a(h[14]) );
    inv_1 \U14/Uil  ( .x(\U14/nl ), .a(l[14]) );
    ao23_1 \U14/Ucl/U1/U1  ( .x(l[14]), .a(n6), .b(l[14]), .c(n1), .d(\U14/ni 
        ), .e(\U14/nh ) );
    ao23_1 \U14/Uch/U1/U1  ( .x(h[14]), .a(n6), .b(h[14]), .c(n3), .d(i[14]), 
        .e(\U14/nl ) );
    inv_1 \U13/Uii  ( .x(\U13/ni ), .a(i[13]) );
    inv_1 \U13/Uih  ( .x(\U13/nh ), .a(h[13]) );
    inv_1 \U13/Uil  ( .x(\U13/nl ), .a(l[13]) );
    ao23_1 \U13/Ucl/U1/U1  ( .x(l[13]), .a(n6), .b(l[13]), .c(n4), .d(\U13/ni 
        ), .e(\U13/nh ) );
    ao23_1 \U13/Uch/U1/U1  ( .x(h[13]), .a(n6), .b(h[13]), .c(n4), .d(i[13]), 
        .e(\U13/nl ) );
    inv_1 \U12/Uii  ( .x(\U12/ni ), .a(i[12]) );
    inv_1 \U12/Uih  ( .x(\U12/nh ), .a(h[12]) );
    inv_1 \U12/Uil  ( .x(\U12/nl ), .a(l[12]) );
    ao23_1 \U12/Ucl/U1/U1  ( .x(l[12]), .a(n5), .b(l[12]), .c(n4), .d(\U12/ni 
        ), .e(\U12/nh ) );
    ao23_1 \U12/Uch/U1/U1  ( .x(h[12]), .a(n5), .b(h[12]), .c(n4), .d(i[12]), 
        .e(\U12/nl ) );
    inv_1 \U11/Uii  ( .x(\U11/ni ), .a(i[11]) );
    inv_1 \U11/Uih  ( .x(\U11/nh ), .a(h[11]) );
    inv_1 \U11/Uil  ( .x(\U11/nl ), .a(l[11]) );
    ao23_1 \U11/Ucl/U1/U1  ( .x(l[11]), .a(n5), .b(l[11]), .c(n4), .d(\U11/ni 
        ), .e(\U11/nh ) );
    ao23_1 \U11/Uch/U1/U1  ( .x(h[11]), .a(n5), .b(h[11]), .c(n4), .d(i[11]), 
        .e(\U11/nl ) );
    inv_1 \U10/Uii  ( .x(\U10/ni ), .a(i[10]) );
    inv_1 \U10/Uih  ( .x(\U10/nh ), .a(h[10]) );
    inv_1 \U10/Uil  ( .x(\U10/nl ), .a(l[10]) );
    ao23_1 \U10/Ucl/U1/U1  ( .x(l[10]), .a(n5), .b(l[10]), .c(n3), .d(\U10/ni 
        ), .e(\U10/nh ) );
    ao23_1 \U10/Uch/U1/U1  ( .x(h[10]), .a(n5), .b(h[10]), .c(n3), .d(i[10]), 
        .e(\U10/nl ) );
    inv_1 \U9/Uii  ( .x(\U9/ni ), .a(i[9]) );
    inv_1 \U9/Uih  ( .x(\U9/nh ), .a(h[9]) );
    inv_1 \U9/Uil  ( .x(\U9/nl ), .a(l[9]) );
    ao23_1 \U9/Ucl/U1/U1  ( .x(l[9]), .a(n5), .b(l[9]), .c(n3), .d(\U9/ni ), 
        .e(\U9/nh ) );
    ao23_1 \U9/Uch/U1/U1  ( .x(h[9]), .a(n5), .b(h[9]), .c(n3), .d(i[9]), .e(
        \U9/nl ) );
    inv_1 \U8/Uii  ( .x(\U8/ni ), .a(i[8]) );
    inv_1 \U8/Uih  ( .x(\U8/nh ), .a(h[8]) );
    inv_1 \U8/Uil  ( .x(\U8/nl ), .a(l[8]) );
    ao23_1 \U8/Ucl/U1/U1  ( .x(l[8]), .a(n5), .b(l[8]), .c(n3), .d(\U8/ni ), 
        .e(\U8/nh ) );
    ao23_1 \U8/Uch/U1/U1  ( .x(h[8]), .a(n5), .b(h[8]), .c(n3), .d(i[8]), .e(
        \U8/nl ) );
    inv_1 \U7/Uii  ( .x(\U7/ni ), .a(i[7]) );
    inv_1 \U7/Uih  ( .x(\U7/nh ), .a(h[7]) );
    inv_1 \U7/Uil  ( .x(\U7/nl ), .a(l[7]) );
    ao23_1 \U7/Ucl/U1/U1  ( .x(l[7]), .a(n7), .b(l[7]), .c(n3), .d(\U7/ni ), 
        .e(\U7/nh ) );
    ao23_1 \U7/Uch/U1/U1  ( .x(h[7]), .a(n7), .b(h[7]), .c(n2), .d(i[7]), .e(
        \U7/nl ) );
    inv_1 \U6/Uii  ( .x(\U6/ni ), .a(i[6]) );
    inv_1 \U6/Uih  ( .x(\U6/nh ), .a(h[6]) );
    inv_1 \U6/Uil  ( .x(\U6/nl ), .a(l[6]) );
    ao23_1 \U6/Ucl/U1/U1  ( .x(l[6]), .a(n7), .b(l[6]), .c(n2), .d(\U6/ni ), 
        .e(\U6/nh ) );
    ao23_1 \U6/Uch/U1/U1  ( .x(h[6]), .a(n7), .b(h[6]), .c(n2), .d(i[6]), .e(
        \U6/nl ) );
    inv_1 \U5/Uii  ( .x(\U5/ni ), .a(i[5]) );
    inv_1 \U5/Uih  ( .x(\U5/nh ), .a(h[5]) );
    inv_1 \U5/Uil  ( .x(\U5/nl ), .a(l[5]) );
    ao23_1 \U5/Ucl/U1/U1  ( .x(l[5]), .a(n7), .b(l[5]), .c(n2), .d(\U5/ni ), 
        .e(\U5/nh ) );
    ao23_1 \U5/Uch/U1/U1  ( .x(h[5]), .a(n7), .b(h[5]), .c(n2), .d(i[5]), .e(
        \U5/nl ) );
    inv_1 \U4/Uii  ( .x(\U4/ni ), .a(i[4]) );
    inv_1 \U4/Uih  ( .x(\U4/nh ), .a(h[4]) );
    inv_1 \U4/Uil  ( .x(\U4/nl ), .a(l[4]) );
    ao23_1 \U4/Ucl/U1/U1  ( .x(l[4]), .a(n6), .b(l[4]), .c(n2), .d(\U4/ni ), 
        .e(\U4/nh ) );
    ao23_1 \U4/Uch/U1/U1  ( .x(h[4]), .a(n6), .b(h[4]), .c(n2), .d(i[4]), .e(
        \U4/nl ) );
    inv_1 \U3/Uii  ( .x(\U3/ni ), .a(i[3]) );
    inv_1 \U3/Uih  ( .x(\U3/nh ), .a(h[3]) );
    inv_1 \U3/Uil  ( .x(\U3/nl ), .a(l[3]) );
    ao23_1 \U3/Ucl/U1/U1  ( .x(l[3]), .a(n6), .b(l[3]), .c(n2), .d(\U3/ni ), 
        .e(\U3/nh ) );
    ao23_1 \U3/Uch/U1/U1  ( .x(h[3]), .a(n8), .b(h[3]), .c(n1), .d(i[3]), .e(
        \U3/nl ) );
    inv_1 \U2/Uii  ( .x(\U2/ni ), .a(i[2]) );
    inv_1 \U2/Uih  ( .x(\U2/nh ), .a(h[2]) );
    inv_1 \U2/Uil  ( .x(\U2/nl ), .a(l[2]) );
    ao23_1 \U2/Ucl/U1/U1  ( .x(l[2]), .a(n8), .b(l[2]), .c(n1), .d(\U2/ni ), 
        .e(\U2/nh ) );
    ao23_1 \U2/Uch/U1/U1  ( .x(h[2]), .a(n8), .b(h[2]), .c(n1), .d(i[2]), .e(
        \U2/nl ) );
    inv_1 \U1/Uii  ( .x(\U1/ni ), .a(i[1]) );
    inv_1 \U1/Uih  ( .x(\U1/nh ), .a(h[1]) );
    inv_1 \U1/Uil  ( .x(\U1/nl ), .a(l[1]) );
    ao23_1 \U1/Ucl/U1/U1  ( .x(l[1]), .a(n8), .b(l[1]), .c(n1), .d(\U1/ni ), 
        .e(\U1/nh ) );
    ao23_1 \U1/Uch/U1/U1  ( .x(h[1]), .a(n8), .b(h[1]), .c(n1), .d(i[1]), .e(
        \U1/nl ) );
    inv_1 \U0/Uii  ( .x(\U0/ni ), .a(i[0]) );
    inv_1 \U0/Uih  ( .x(\U0/nh ), .a(h[0]) );
    inv_1 \U0/Uil  ( .x(\U0/nl ), .a(l[0]) );
    ao23_1 \U0/Ucl/U1/U1  ( .x(l[0]), .a(n8), .b(l[0]), .c(n1), .d(\U0/ni ), 
        .e(\U0/nh ) );
    ao23_1 \U0/Uch/U1/U1  ( .x(h[0]), .a(n8), .b(h[0]), .c(n1), .d(i[0]), .e(
        \U0/nl ) );
    buf_16 U1 ( .x(n1), .a(n12) );
    buf_16 U2 ( .x(n2), .a(n12) );
    buf_16 U3 ( .x(n3), .a(n12) );
    buf_16 U4 ( .x(n4), .a(n11) );
    buf_16 U5 ( .x(n5), .a(n11) );
    buf_16 U6 ( .x(n6), .a(n11) );
    buf_16 U7 ( .x(n7), .a(n10) );
    buf_16 U8 ( .x(n8), .a(n10) );
    buf_16 U9 ( .x(n9), .a(n10) );
    buf_16 U10 ( .x(n10), .a(req) );
    buf_16 U11 ( .x(n11), .a(req) );
    buf_16 U12 ( .x(n12), .a(req) );
endmodule


module latch_ctrl_2 ( rin, ain, rout, aout, en, reset );
input  rin, aout, reset;
output ain, rout, en;
    wire N5, N6, na, a, n_rout, nreset, n3, \c_rout/ob , n1;
    inv_1 U0 ( .x(nreset), .a(reset) );
    nor2_1 U1 ( .x(ain), .a(na), .b(n1) );
    inv_1 U2 ( .x(na), .a(a) );
    inv_1 U3 ( .x(N6), .a(N5) );
    and2_1 C9 ( .x(n3), .a(na), .b(N6) );
    or2_1 C11 ( .x(N5), .a(rout), .b(aout) );
    oa21_1 \c_na/__tmp99/U1  ( .x(a), .a(n1), .b(a), .c(rin) );
    oai21_1 \c_rout/U1  ( .x(\c_rout/ob ), .a(aout), .b(n_rout), .c(na) );
    nand2_1 \c_rout/U2  ( .x(n_rout), .a(nreset), .b(\c_rout/ob ) );
    buf_1 U4 ( .x(en), .a(n3) );
    inv_2 U5 ( .x(rout), .a(n_rout) );
    buf_1 U6 ( .x(n1), .a(n3) );
endmodule


module m2cp_tic ( req_in, ts_o, sel_o, mult_o, we_o, prd_o, seq_o, adr_o, 
    dat_o, ain, ic_seq, ic_pred, ic_size, ic_itag, ic_wd, ic_lock, ic_a, 
    ic_rnw, ic_col, ic_ack, req_out, ts_i, we_i, err_i, rty_i, acc_i, dat_i, 
    aout, ir_rd, ir_err, ir_rnw, ir_ack, tag_id, reset );
input  [2:0] ts_o;
input  [3:0] sel_o;
input  [31:0] adr_o;
input  [31:0] dat_o;
output [1:0] ic_seq;
output [1:0] ic_pred;
output [3:0] ic_size;
output [9:0] ic_itag;
output [63:0] ic_wd;
output [1:0] ic_lock;
output [63:0] ic_a;
output [1:0] ic_rnw;
output [5:0] ic_col;
output [2:0] ts_i;
output [31:0] dat_i;
input  [63:0] ir_rd;
input  [1:0] ir_err;
input  [1:0] ir_rnw;
input  [4:0] tag_id;
input  req_in, mult_o, we_o, prd_o, seq_o, ic_ack, aout, reset;
output ain, req_out, we_i, err_i, rty_i, acc_i, ir_ack;
    wire n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
        n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, 
        n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, 
        n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
        n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
        n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
        n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
        n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
        n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
        n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
        n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
        n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
        n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
        n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
        n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
        n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
        n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
        n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
        n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
        n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
        n308, n2, n3, n4, n5, req_in_delayed, \size[1] , \size[0] , \data[15] , 
        \data[14] , \data[13] , \data[12] , \data[11] , \data[10] , \data[9] , 
        \data[8] , \data[7] , \data[6] , \data[5] , \data[4] , \data[3] , 
        \data[2] , \data[1] , \data[0] , _24_net_, _25_net_, _26_net_, 
        comp_basic, high_ir_rd, low_ir_rd, comp_rd, _27_net_, all_r, _28_net_, 
        all_w, complete, complete_delayed, en, \all_read/__tmp99/loop , 
        \Ucol2/nl , \Ucol2/ni , \Ucol2/nh , \Ucol1/nl , \Ucol1/ni , \Ucol1/nh , 
        \Ucol0/nl , \Ucol0/ni , \Ucol0/nh , \Utag4/nl , \Utag4/ni , \Utag4/nh , 
        \Utag3/nl , \Utag3/ni , \Utag3/nh , \Utag2/nl , \Utag2/ni , \Utag2/nh , 
        \Utag1/nl , \Utag1/ni , \Utag1/nh , \Utag0/nl , \Utag0/ni , \Utag0/nh , 
        \Usze1/nl , \Usze1/ni , \Usze1/nh , \Usze0/nl , \Usze0/ni , \Usze0/nh , 
        \Urnw/nl , \Urnw/ni , \Urnw/nh , \Ulock/nl , \Ulock/ni , \Ulock/nh , 
        \Upred/nl , \Upred/ni , \Upred/nh , \Useq/nl , \Useq/ni , \Useq/nh , 
        n1, n6, n7, n8, n9, n10, n11;
    assign ain = ic_ack;
    assign ts_i[2] = 1'b0;
    assign ts_i[1] = 1'b0;
    assign ts_i[0] = 1'b0;
    assign rty_i = 1'b0;
    assign acc_i = 1'b0;
    matched_delay_m2cp_com_tic U130 ( .x(req_in_delayed), .a(req_in) );
    sr2dr_word_5 Uwd ( .i({dat_o[31], dat_o[30], dat_o[29], dat_o[28], 
        dat_o[27], dat_o[26], dat_o[25], dat_o[24], dat_o[23], dat_o[22], 
        dat_o[21], dat_o[20], dat_o[19], dat_o[18], dat_o[17], dat_o[16], 
        \data[15] , \data[14] , \data[13] , \data[12] , \data[11] , \data[10] , 
        \data[9] , \data[8] , \data[7] , \data[6] , \data[5] , \data[4] , 
        \data[3] , \data[2] , \data[1] , \data[0] }), .req(n8), .h(ic_wd
        [63:32]), .l(ic_wd[31:0]) );
    sr2dr_word_4 Ua ( .i(adr_o), .req(n8), .h(ic_a[63:32]), .l(ic_a[31:0]) );
    latch_ctrl_2 lc ( .rin(complete_delayed), .ain(ir_ack), .rout(req_out), 
        .aout(aout), .en(en), .reset(reset) );
    nand2_1 U61 ( .x(_26_net_), .a(n72), .b(n77) );
    and2_1 U274 ( .x(_27_net_), .a(ir_rnw[1]), .b(ir_err[0]) );
    inv_1 U275 ( .x(_24_net_), .a(we_o) );
    inv_1 U2 ( .x(n112), .a(ir_rd[4]) );
    inv_1 U3 ( .x(n124), .a(ir_rd[0]) );
    inv_1 U4 ( .x(n118), .a(ir_rd[2]) );
    inv_1 U5 ( .x(n206), .a(dat_o[28]) );
    inv_1 U6 ( .x(n208), .a(dat_o[27]) );
    inv_1 U7 ( .x(n210), .a(dat_o[26]) );
    inv_1 U8 ( .x(n197), .a(dat_o[25]) );
    inv_1 U9 ( .x(n199), .a(dat_o[24]) );
    inv_1 U10 ( .x(n202), .a(dat_o[15]) );
    inv_1 U11 ( .x(n201), .a(dat_o[31]) );
    inv_1 U12 ( .x(n203), .a(dat_o[30]) );
    inv_1 U13 ( .x(n204), .a(dat_o[29]) );
    nor2_1 U14 ( .x(\size[1] ), .a(n83), .b(n84) );
    inv_1 U15 ( .x(n72), .a(ir_rnw[0]) );
    oa21_1 U16 ( .x(n89), .a(n205), .b(n64), .c(n2) );
    inv_1 U24 ( .x(n2), .a(n90) );
    inv_1 U17 ( .x(n205), .a(dat_o[13]) );
    inv_1 U18 ( .x(n64), .a(sel_o[1]) );
    oa21_1 U19 ( .x(n97), .a(n198), .b(n64), .c(n3) );
    inv_1 U276 ( .x(n3), .a(n98) );
    inv_1 U20 ( .x(n198), .a(dat_o[9]) );
    oa21_1 U21 ( .x(n87), .a(n63), .b(n64), .c(n4) );
    inv_1 U277 ( .x(n4), .a(n88) );
    inv_1 U22 ( .x(n63), .a(dat_o[14]) );
    oa21_1 U23 ( .x(n85), .a(n202), .b(n64), .c(n5) );
    inv_1 U278 ( .x(n5), .a(n86) );
    nand2_1 U25 ( .x(n290), .a(n289), .b(n288) );
    nand2_1 U26 ( .x(n79), .a(n277), .b(n270) );
    nor2_1 U27 ( .x(n277), .a(n273), .b(n276) );
    nor2_1 U28 ( .x(n270), .a(n266), .b(n269) );
    nand2_1 U29 ( .x(n283), .a(n282), .b(n281) );
    nand2_1 U30 ( .x(n298), .a(dat_o[20]), .b(n70) );
    inv_1 U31 ( .x(n70), .a(n68) );
    nand2_1 U32 ( .x(n213), .a(n223), .b(n71) );
    nand2_1 U33 ( .x(n80), .a(n291), .b(n284) );
    nor2_1 U34 ( .x(n291), .a(n287), .b(n290) );
    nor2_1 U35 ( .x(n284), .a(n280), .b(n283) );
    aoi21_1 U36 ( .x(n99), .a(dat_o[8]), .b(n71), .c(n100) );
    aoi21_1 U37 ( .x(n95), .a(dat_o[10]), .b(n71), .c(n96) );
    aoi21_1 U38 ( .x(n93), .a(dat_o[11]), .b(n71), .c(n94) );
    aoi21_1 U39 ( .x(n91), .a(dat_o[12]), .b(n71), .c(n92) );
    inv_1 U40 ( .x(n81), .a(all_r) );
    buf_1 U41 ( .x(n65), .a(sel_o[0]) );
    nand2_1 U42 ( .x(n84), .a(sel_o[0]), .b(n71) );
    inv_1 U43 ( .x(n66), .a(sel_o[3]) );
    inv_1 U44 ( .x(n67), .a(n66) );
    inv_1 U45 ( .x(n68), .a(sel_o[2]) );
    inv_1 U46 ( .x(n69), .a(n68) );
    nand2_1 U48 ( .x(n83), .a(n70), .b(n67) );
    nand3i_1 U49 ( .x(n212), .a(sel_o[1]), .b(n67), .c(n70) );
    nor2_1 U50 ( .x(n223), .a(n70), .b(n67) );
    nand2_1 U51 ( .x(n300), .a(dat_o[19]), .b(n69) );
    nand2_1 U52 ( .x(n294), .a(dat_o[22]), .b(n69) );
    nand2_1 U53 ( .x(n302), .a(dat_o[18]), .b(n69) );
    nand2_1 U54 ( .x(n296), .a(dat_o[21]), .b(n69) );
    nand2_1 U55 ( .x(n306), .a(dat_o[16]), .b(n69) );
    nand2_1 U56 ( .x(n292), .a(dat_o[23]), .b(n69) );
    nand2_1 U57 ( .x(n304), .a(dat_o[17]), .b(n69) );
    buf_1 U58 ( .x(n71), .a(sel_o[1]) );
    nand4_1 U60 ( .x(low_ir_rd), .a(n73), .b(n74), .c(n75), .d(n76) );
    nand2_1 U62 ( .x(complete), .a(n81), .b(n82) );
    matched_delay_m2cp_resp_tic mdel ( .x(complete_delayed), .a(complete) );
    inv_1 U63 ( .x(n200), .a(dat_o[8]) );
    inv_1 U64 ( .x(n207), .a(dat_o[12]) );
    inv_1 U65 ( .x(n209), .a(dat_o[11]) );
    inv_1 U66 ( .x(n211), .a(dat_o[10]) );
    nand4_1 U67 ( .x(n224), .a(n225), .b(n226), .c(n227), .d(n228) );
    nand4_1 U68 ( .x(n229), .a(n230), .b(n231), .c(n232), .d(n233) );
    nor2_1 U69 ( .x(n76), .a(n224), .b(n229) );
    nand4_1 U70 ( .x(n234), .a(n235), .b(n236), .c(n237), .d(n238) );
    nand4_1 U71 ( .x(n239), .a(n240), .b(n241), .c(n242), .d(n243) );
    nor2_1 U72 ( .x(n75), .a(n234), .b(n239) );
    nand4_1 U73 ( .x(n244), .a(n245), .b(n246), .c(n247), .d(n248) );
    nand4_1 U74 ( .x(n249), .a(n250), .b(n251), .c(n252), .d(n253) );
    nor2_1 U75 ( .x(n74), .a(n244), .b(n249) );
    nand4_1 U76 ( .x(n254), .a(n255), .b(n256), .c(n257), .d(n258) );
    nand4_1 U77 ( .x(n259), .a(n260), .b(n261), .c(n262), .d(n263) );
    nor2_1 U78 ( .x(n73), .a(n254), .b(n259) );
    nand2_1 U79 ( .x(n266), .a(n265), .b(n264) );
    nand2_1 U80 ( .x(n269), .a(n268), .b(n267) );
    nand2_1 U81 ( .x(n273), .a(n272), .b(n271) );
    nand2_1 U82 ( .x(n276), .a(n275), .b(n274) );
    nand2_1 U83 ( .x(n280), .a(n279), .b(n278) );
    nand2_1 U84 ( .x(n287), .a(n286), .b(n285) );
    nand2_1 U85 ( .x(n86), .a(n292), .b(n293) );
    nand2_1 U86 ( .x(n88), .a(n294), .b(n295) );
    nand2_1 U87 ( .x(n90), .a(n296), .b(n297) );
    nand2_1 U88 ( .x(n92), .a(n298), .b(n299) );
    nand2_1 U89 ( .x(n94), .a(n300), .b(n301) );
    nand2_1 U90 ( .x(n96), .a(n302), .b(n303) );
    nand2_1 U91 ( .x(n98), .a(n304), .b(n305) );
    nand2_1 U92 ( .x(n100), .a(n306), .b(n307) );
    inv_1 U93 ( .x(n222), .a(dat_o[0]) );
    inv_1 U94 ( .x(n221), .a(dat_o[1]) );
    inv_1 U95 ( .x(n220), .a(dat_o[2]) );
    inv_1 U96 ( .x(n219), .a(dat_o[3]) );
    inv_1 U97 ( .x(n218), .a(dat_o[4]) );
    inv_1 U98 ( .x(n217), .a(dat_o[5]) );
    inv_1 U99 ( .x(n216), .a(dat_o[6]) );
    inv_1 U100 ( .x(n215), .a(dat_o[7]) );
    inv_1 U101 ( .x(n77), .a(ir_rnw[1]) );
    inv_1 U103 ( .x(n82), .a(all_w) );
    nand2_1 U104 ( .x(n293), .a(dat_o[31]), .b(n67) );
    nand2_1 U105 ( .x(n295), .a(dat_o[30]), .b(n67) );
    nand2_1 U106 ( .x(n297), .a(dat_o[29]), .b(n67) );
    nand2_1 U107 ( .x(n299), .a(dat_o[28]), .b(n67) );
    nand2_1 U108 ( .x(n301), .a(dat_o[27]), .b(n67) );
    nand2_1 U109 ( .x(n303), .a(dat_o[26]), .b(n67) );
    nand2_1 U110 ( .x(n305), .a(dat_o[25]), .b(n67) );
    nand2_1 U111 ( .x(n307), .a(dat_o[24]), .b(n67) );
    mux2i_1 U113 ( .x(\data[0] ), .d0(n99), .sl(n65), .d1(n222) );
    mux2i_1 U114 ( .x(\data[10] ), .d0(n211), .sl(n214), .d1(n210) );
    mux2i_1 U115 ( .x(\data[11] ), .d0(n209), .sl(n214), .d1(n208) );
    mux2i_1 U116 ( .x(\data[12] ), .d0(n207), .sl(n214), .d1(n206) );
    mux2i_1 U117 ( .x(\data[13] ), .d0(n205), .sl(n214), .d1(n204) );
    mux2i_1 U118 ( .x(\data[14] ), .d0(n63), .sl(n214), .d1(n203) );
    mux2i_1 U119 ( .x(\data[15] ), .d0(n202), .sl(n214), .d1(n201) );
    mux2i_1 U120 ( .x(\data[1] ), .d0(n97), .sl(n65), .d1(n221) );
    mux2i_1 U121 ( .x(\data[2] ), .d0(n95), .sl(n65), .d1(n220) );
    mux2i_1 U122 ( .x(\data[3] ), .d0(n93), .sl(n65), .d1(n219) );
    mux2i_1 U123 ( .x(\data[4] ), .d0(n91), .sl(n65), .d1(n218) );
    mux2i_1 U124 ( .x(\data[5] ), .d0(n89), .sl(n65), .d1(n217) );
    mux2i_1 U125 ( .x(\data[6] ), .d0(n87), .sl(n65), .d1(n216) );
    mux2i_1 U126 ( .x(\data[7] ), .d0(n85), .sl(n65), .d1(n215) );
    mux2i_1 U127 ( .x(\data[8] ), .d0(n200), .sl(n214), .d1(n199) );
    mux2i_1 U128 ( .x(\data[9] ), .d0(n198), .sl(n214), .d1(n197) );
    nor2_1 U129 ( .x(high_ir_rd), .a(n79), .b(n80) );
    mux2i_1 U131 ( .x(\size[0] ), .d0(n212), .sl(n65), .d1(n213) );
    nand2i_1 U132 ( .x(n308), .a(sel_o[1]), .b(n70) );
    inv_1 U133 ( .x(n255), .a(n182) );
    inv_1 U134 ( .x(n256), .a(n179) );
    inv_1 U135 ( .x(n257), .a(n176) );
    inv_1 U136 ( .x(n258), .a(n173) );
    inv_1 U137 ( .x(n260), .a(n194) );
    inv_1 U138 ( .x(n261), .a(n191) );
    inv_1 U139 ( .x(n262), .a(n188) );
    inv_1 U140 ( .x(n263), .a(n185) );
    inv_1 U141 ( .x(n245), .a(n158) );
    inv_1 U142 ( .x(n246), .a(n155) );
    inv_1 U143 ( .x(n247), .a(n152) );
    inv_1 U144 ( .x(n248), .a(n149) );
    inv_1 U145 ( .x(n250), .a(n170) );
    inv_1 U146 ( .x(n251), .a(n167) );
    inv_1 U147 ( .x(n252), .a(n164) );
    inv_1 U148 ( .x(n253), .a(n161) );
    inv_1 U149 ( .x(n235), .a(n134) );
    inv_1 U150 ( .x(n236), .a(n131) );
    inv_1 U151 ( .x(n237), .a(n128) );
    inv_1 U152 ( .x(n238), .a(n125) );
    inv_1 U153 ( .x(n240), .a(n146) );
    inv_1 U154 ( .x(n241), .a(n143) );
    inv_1 U155 ( .x(n242), .a(n140) );
    inv_1 U156 ( .x(n243), .a(n137) );
    inv_1 U157 ( .x(n225), .a(n110) );
    inv_1 U158 ( .x(n226), .a(n107) );
    inv_1 U159 ( .x(n227), .a(n104) );
    inv_1 U160 ( .x(n228), .a(n101) );
    inv_1 U161 ( .x(n230), .a(n122) );
    inv_1 U162 ( .x(n231), .a(n119) );
    inv_1 U163 ( .x(n232), .a(n116) );
    inv_1 U164 ( .x(n233), .a(n113) );
    nor2_1 U165 ( .x(n272), .a(n252), .b(n253) );
    nor2_1 U166 ( .x(n271), .a(n250), .b(n251) );
    nor2_1 U167 ( .x(n275), .a(n247), .b(n248) );
    nor2_1 U168 ( .x(n274), .a(n245), .b(n246) );
    nor2_1 U169 ( .x(n265), .a(n262), .b(n263) );
    nor2_1 U170 ( .x(n264), .a(n260), .b(n261) );
    nor2_1 U171 ( .x(n268), .a(n257), .b(n258) );
    nor2_1 U172 ( .x(n267), .a(n255), .b(n256) );
    nor2_1 U173 ( .x(n286), .a(n232), .b(n233) );
    nor2_1 U174 ( .x(n285), .a(n230), .b(n231) );
    nor2_1 U175 ( .x(n289), .a(n227), .b(n228) );
    nor2_1 U176 ( .x(n288), .a(n225), .b(n226) );
    nor2_1 U177 ( .x(n279), .a(n242), .b(n243) );
    nor2_1 U178 ( .x(n278), .a(n240), .b(n241) );
    nor2_1 U179 ( .x(n282), .a(n237), .b(n238) );
    nor2_1 U180 ( .x(n281), .a(n235), .b(n236) );
    nand2_1 U181 ( .x(n182), .a(n183), .b(n184) );
    nand2_1 U182 ( .x(n179), .a(n180), .b(n181) );
    nand2_1 U183 ( .x(n176), .a(n177), .b(n178) );
    nand2_1 U184 ( .x(n173), .a(n174), .b(n175) );
    nand2_1 U185 ( .x(n194), .a(n195), .b(n196) );
    nand2_1 U186 ( .x(n191), .a(n192), .b(n193) );
    nand2_1 U187 ( .x(n188), .a(n189), .b(n190) );
    nand2_1 U188 ( .x(n185), .a(n186), .b(n187) );
    nand2_1 U189 ( .x(n158), .a(n159), .b(n160) );
    nand2_1 U190 ( .x(n155), .a(n156), .b(n157) );
    nand2_1 U191 ( .x(n152), .a(n153), .b(n154) );
    nand2_1 U192 ( .x(n149), .a(n150), .b(n151) );
    nand2_1 U193 ( .x(n170), .a(n171), .b(n172) );
    nand2_1 U194 ( .x(n167), .a(n168), .b(n169) );
    nand2_1 U195 ( .x(n164), .a(n165), .b(n166) );
    nand2_1 U196 ( .x(n161), .a(n162), .b(n163) );
    nand2_1 U197 ( .x(n134), .a(n135), .b(n136) );
    nand2_1 U198 ( .x(n131), .a(n132), .b(n133) );
    nand2_1 U199 ( .x(n128), .a(n129), .b(n130) );
    nand2_1 U200 ( .x(n125), .a(n126), .b(n127) );
    nand2_1 U201 ( .x(n146), .a(n147), .b(n148) );
    nand2_1 U202 ( .x(n143), .a(n144), .b(n145) );
    nand2_1 U203 ( .x(n140), .a(n141), .b(n142) );
    nand2_1 U204 ( .x(n137), .a(n138), .b(n139) );
    nand2_1 U205 ( .x(n110), .a(n111), .b(n112) );
    nand2_1 U206 ( .x(n107), .a(n108), .b(n109) );
    nand2_1 U207 ( .x(n104), .a(n105), .b(n106) );
    nand2_1 U208 ( .x(n101), .a(n102), .b(n103) );
    nand2_1 U209 ( .x(n122), .a(n123), .b(n124) );
    nand2_1 U210 ( .x(n119), .a(n120), .b(n121) );
    nand2_1 U211 ( .x(n116), .a(n117), .b(n118) );
    nand2_1 U212 ( .x(n113), .a(n114), .b(n115) );
    inv_1 U213 ( .x(n183), .a(ir_rd[60]) );
    inv_1 U214 ( .x(n184), .a(ir_rd[28]) );
    inv_1 U215 ( .x(n180), .a(ir_rd[61]) );
    inv_1 U216 ( .x(n181), .a(ir_rd[29]) );
    inv_1 U217 ( .x(n177), .a(ir_rd[62]) );
    inv_1 U218 ( .x(n178), .a(ir_rd[30]) );
    inv_1 U219 ( .x(n174), .a(ir_rd[63]) );
    inv_1 U220 ( .x(n175), .a(ir_rd[31]) );
    inv_1 U221 ( .x(n195), .a(ir_rd[56]) );
    inv_1 U222 ( .x(n196), .a(ir_rd[24]) );
    inv_1 U223 ( .x(n192), .a(ir_rd[57]) );
    inv_1 U224 ( .x(n193), .a(ir_rd[25]) );
    inv_1 U225 ( .x(n189), .a(ir_rd[58]) );
    inv_1 U226 ( .x(n190), .a(ir_rd[26]) );
    inv_1 U227 ( .x(n186), .a(ir_rd[59]) );
    inv_1 U228 ( .x(n187), .a(ir_rd[27]) );
    inv_1 U229 ( .x(n159), .a(ir_rd[52]) );
    inv_1 U230 ( .x(n160), .a(ir_rd[20]) );
    inv_1 U231 ( .x(n156), .a(ir_rd[53]) );
    inv_1 U232 ( .x(n157), .a(ir_rd[21]) );
    inv_1 U233 ( .x(n153), .a(ir_rd[54]) );
    inv_1 U234 ( .x(n154), .a(ir_rd[22]) );
    inv_1 U235 ( .x(n150), .a(ir_rd[55]) );
    inv_1 U236 ( .x(n151), .a(ir_rd[23]) );
    inv_1 U237 ( .x(n171), .a(ir_rd[48]) );
    inv_1 U238 ( .x(n172), .a(ir_rd[16]) );
    inv_1 U239 ( .x(n168), .a(ir_rd[49]) );
    inv_1 U240 ( .x(n169), .a(ir_rd[17]) );
    inv_1 U241 ( .x(n165), .a(ir_rd[50]) );
    inv_1 U242 ( .x(n166), .a(ir_rd[18]) );
    inv_1 U243 ( .x(n162), .a(ir_rd[51]) );
    inv_1 U244 ( .x(n163), .a(ir_rd[19]) );
    inv_1 U245 ( .x(n135), .a(ir_rd[44]) );
    inv_1 U246 ( .x(n136), .a(ir_rd[12]) );
    inv_1 U247 ( .x(n132), .a(ir_rd[45]) );
    inv_1 U248 ( .x(n133), .a(ir_rd[13]) );
    inv_1 U249 ( .x(n129), .a(ir_rd[46]) );
    inv_1 U250 ( .x(n130), .a(ir_rd[14]) );
    inv_1 U251 ( .x(n126), .a(ir_rd[47]) );
    inv_1 U252 ( .x(n127), .a(ir_rd[15]) );
    inv_1 U253 ( .x(n147), .a(ir_rd[40]) );
    inv_1 U254 ( .x(n148), .a(ir_rd[8]) );
    inv_1 U255 ( .x(n144), .a(ir_rd[41]) );
    inv_1 U256 ( .x(n145), .a(ir_rd[9]) );
    inv_1 U257 ( .x(n141), .a(ir_rd[42]) );
    inv_1 U258 ( .x(n142), .a(ir_rd[10]) );
    inv_1 U259 ( .x(n138), .a(ir_rd[43]) );
    inv_1 U260 ( .x(n139), .a(ir_rd[11]) );
    inv_1 U261 ( .x(n111), .a(ir_rd[36]) );
    inv_1 U262 ( .x(n108), .a(ir_rd[37]) );
    inv_1 U263 ( .x(n109), .a(ir_rd[5]) );
    inv_1 U264 ( .x(n105), .a(ir_rd[38]) );
    inv_1 U265 ( .x(n106), .a(ir_rd[6]) );
    inv_1 U266 ( .x(n102), .a(ir_rd[39]) );
    inv_1 U267 ( .x(n103), .a(ir_rd[7]) );
    inv_1 U268 ( .x(n123), .a(ir_rd[32]) );
    inv_1 U269 ( .x(n120), .a(ir_rd[33]) );
    inv_1 U270 ( .x(n121), .a(ir_rd[1]) );
    inv_1 U271 ( .x(n117), .a(ir_rd[34]) );
    inv_1 U272 ( .x(n114), .a(ir_rd[35]) );
    inv_1 U273 ( .x(n115), .a(ir_rd[3]) );
    latn_1 \dat_i_reg[30]  ( .q(dat_i[30]), .d(ir_rd[62]), .g(n7) );
    latn_1 \dat_i_reg[28]  ( .q(dat_i[28]), .d(ir_rd[60]), .g(n7) );
    latn_1 \dat_i_reg[27]  ( .q(dat_i[27]), .d(ir_rd[59]), .g(n7) );
    latn_1 \dat_i_reg[26]  ( .q(dat_i[26]), .d(ir_rd[58]), .g(n7) );
    latn_1 \dat_i_reg[25]  ( .q(dat_i[25]), .d(ir_rd[57]), .g(n7) );
    latn_1 \dat_i_reg[24]  ( .q(dat_i[24]), .d(ir_rd[56]), .g(n7) );
    latn_1 \dat_i_reg[22]  ( .q(dat_i[22]), .d(ir_rd[54]), .g(n7) );
    latn_1 \dat_i_reg[20]  ( .q(dat_i[20]), .d(ir_rd[52]), .g(n7) );
    latn_1 \dat_i_reg[19]  ( .q(dat_i[19]), .d(ir_rd[51]), .g(n7) );
    latn_1 \dat_i_reg[18]  ( .q(dat_i[18]), .d(ir_rd[50]), .g(n7) );
    latn_1 \dat_i_reg[17]  ( .q(dat_i[17]), .d(ir_rd[49]), .g(n7) );
    latn_1 \dat_i_reg[16]  ( .q(dat_i[16]), .d(ir_rd[48]), .g(n6) );
    latn_1 \dat_i_reg[14]  ( .q(dat_i[14]), .d(ir_rd[46]), .g(n6) );
    latn_1 \dat_i_reg[12]  ( .q(dat_i[12]), .d(ir_rd[44]), .g(n6) );
    latn_1 \dat_i_reg[10]  ( .q(dat_i[10]), .d(ir_rd[42]), .g(n6) );
    latn_1 \dat_i_reg[8]  ( .q(dat_i[8]), .d(ir_rd[40]), .g(n6) );
    latn_1 \dat_i_reg[6]  ( .q(dat_i[6]), .d(ir_rd[38]), .g(n6) );
    latn_1 \dat_i_reg[4]  ( .q(dat_i[4]), .d(ir_rd[36]), .g(n6) );
    latn_1 \dat_i_reg[3]  ( .q(dat_i[3]), .d(ir_rd[35]), .g(n1) );
    latn_1 \dat_i_reg[2]  ( .q(dat_i[2]), .d(ir_rd[34]), .g(n1) );
    latn_1 \dat_i_reg[1]  ( .q(dat_i[1]), .d(ir_rd[33]), .g(n1) );
    latn_1 \dat_i_reg[0]  ( .q(dat_i[0]), .d(ir_rd[32]), .g(n1) );
    latn_1 we_i_reg ( .q(we_i), .d(ir_rnw[0]), .g(n1) );
    latn_1 err_i_reg ( .q(err_i), .d(ir_err[1]), .g(n1) );
    latn_1 \dat_i_reg[13]  ( .q(dat_i[13]), .d(ir_rd[45]), .g(n6) );
    latn_1 \dat_i_reg[5]  ( .q(dat_i[5]), .d(ir_rd[37]), .g(n1) );
    latn_1 \dat_i_reg[15]  ( .q(dat_i[15]), .d(ir_rd[47]), .g(n6) );
    latn_1 \dat_i_reg[7]  ( .q(dat_i[7]), .d(ir_rd[39]), .g(n1) );
    latn_1 \dat_i_reg[29]  ( .q(dat_i[29]), .d(ir_rd[61]), .g(n6) );
    latn_1 \dat_i_reg[21]  ( .q(dat_i[21]), .d(ir_rd[53]), .g(n1) );
    latn_1 \dat_i_reg[31]  ( .q(dat_i[31]), .d(ir_rd[63]), .g(n6) );
    latn_1 \dat_i_reg[23]  ( .q(dat_i[23]), .d(ir_rd[55]), .g(n1) );
    latn_1 \dat_i_reg[9]  ( .q(dat_i[9]), .d(ir_rd[41]), .g(n6) );
    latn_1 \dat_i_reg[11]  ( .q(dat_i[11]), .d(ir_rd[43]), .g(n1) );
    oa21_1 \all_write/__tmp99/U1  ( .x(all_w), .a(_28_net_), .b(all_w), .c(
        comp_basic) );
    ao31_1 \all_read/__tmp99/aoi  ( .x(\all_read/__tmp99/loop ), .a(comp_basic
        ), .b(comp_rd), .c(_27_net_), .d(all_r) );
    oa21_1 \all_read/__tmp99/outGate  ( .x(all_r), .a(comp_basic), .b(comp_rd), 
        .c(\all_read/__tmp99/loop ) );
    ao222_1 \rd/__tmp99/U1  ( .x(comp_rd), .a(high_ir_rd), .b(low_ir_rd), .c(
        high_ir_rd), .d(comp_rd), .e(low_ir_rd), .f(comp_rd) );
    ao222_1 \basic/__tmp99/U1  ( .x(comp_basic), .a(_25_net_), .b(_26_net_), 
        .c(_25_net_), .d(comp_basic), .e(_26_net_), .f(comp_basic) );
    inv_1 \Ucol2/Uii  ( .x(\Ucol2/ni ), .a(ts_o[2]) );
    inv_1 \Ucol2/Uih  ( .x(\Ucol2/nh ), .a(ic_col[5]) );
    inv_1 \Ucol2/Uil  ( .x(\Ucol2/nl ), .a(ic_col[2]) );
    ao23_1 \Ucol2/Ucl/U1/U1  ( .x(ic_col[2]), .a(n11), .b(ic_col[2]), .c(n8), 
        .d(\Ucol2/ni ), .e(\Ucol2/nh ) );
    ao23_1 \Ucol2/Uch/U1/U1  ( .x(ic_col[5]), .a(n11), .b(ic_col[5]), .c(n8), 
        .d(ts_o[2]), .e(\Ucol2/nl ) );
    inv_1 \Ucol1/Uii  ( .x(\Ucol1/ni ), .a(ts_o[1]) );
    inv_1 \Ucol1/Uih  ( .x(\Ucol1/nh ), .a(ic_col[4]) );
    inv_1 \Ucol1/Uil  ( .x(\Ucol1/nl ), .a(ic_col[1]) );
    ao23_1 \Ucol1/Ucl/U1/U1  ( .x(ic_col[1]), .a(n11), .b(ic_col[1]), .c(n8), 
        .d(\Ucol1/ni ), .e(\Ucol1/nh ) );
    ao23_1 \Ucol1/Uch/U1/U1  ( .x(ic_col[4]), .a(n11), .b(ic_col[4]), .c(n9), 
        .d(ts_o[1]), .e(\Ucol1/nl ) );
    inv_1 \Ucol0/Uii  ( .x(\Ucol0/ni ), .a(ts_o[0]) );
    inv_1 \Ucol0/Uih  ( .x(\Ucol0/nh ), .a(ic_col[3]) );
    inv_1 \Ucol0/Uil  ( .x(\Ucol0/nl ), .a(ic_col[0]) );
    ao23_1 \Ucol0/Ucl/U1/U1  ( .x(ic_col[0]), .a(n11), .b(ic_col[0]), .c(n10), 
        .d(\Ucol0/ni ), .e(\Ucol0/nh ) );
    ao23_1 \Ucol0/Uch/U1/U1  ( .x(ic_col[3]), .a(n11), .b(ic_col[3]), .c(n9), 
        .d(ts_o[0]), .e(\Ucol0/nl ) );
    inv_1 \Utag4/Uii  ( .x(\Utag4/ni ), .a(tag_id[4]) );
    inv_1 \Utag4/Uih  ( .x(\Utag4/nh ), .a(ic_itag[9]) );
    inv_1 \Utag4/Uil  ( .x(\Utag4/nl ), .a(ic_itag[4]) );
    ao23_1 \Utag4/Ucl/U1/U1  ( .x(ic_itag[4]), .a(n11), .b(ic_itag[4]), .c(n9), 
        .d(\Utag4/ni ), .e(\Utag4/nh ) );
    ao23_1 \Utag4/Uch/U1/U1  ( .x(ic_itag[9]), .a(n10), .b(ic_itag[9]), .c(n9), 
        .d(tag_id[4]), .e(\Utag4/nl ) );
    inv_1 \Utag3/Uii  ( .x(\Utag3/ni ), .a(tag_id[3]) );
    inv_1 \Utag3/Uih  ( .x(\Utag3/nh ), .a(ic_itag[8]) );
    inv_1 \Utag3/Uil  ( .x(\Utag3/nl ), .a(ic_itag[3]) );
    ao23_1 \Utag3/Ucl/U1/U1  ( .x(ic_itag[3]), .a(n10), .b(ic_itag[3]), .c(n9), 
        .d(\Utag3/ni ), .e(\Utag3/nh ) );
    ao23_1 \Utag3/Uch/U1/U1  ( .x(ic_itag[8]), .a(n10), .b(ic_itag[8]), .c(n9), 
        .d(tag_id[3]), .e(\Utag3/nl ) );
    inv_1 \Utag2/Uii  ( .x(\Utag2/ni ), .a(tag_id[2]) );
    inv_1 \Utag2/Uih  ( .x(\Utag2/nh ), .a(ic_itag[7]) );
    inv_1 \Utag2/Uil  ( .x(\Utag2/nl ), .a(ic_itag[2]) );
    ao23_1 \Utag2/Ucl/U1/U1  ( .x(ic_itag[2]), .a(n10), .b(ic_itag[2]), .c(n9), 
        .d(\Utag2/ni ), .e(\Utag2/nh ) );
    ao23_1 \Utag2/Uch/U1/U1  ( .x(ic_itag[7]), .a(n10), .b(ic_itag[7]), .c(n10
        ), .d(tag_id[2]), .e(\Utag2/nl ) );
    inv_1 \Utag1/Uii  ( .x(\Utag1/ni ), .a(tag_id[1]) );
    inv_1 \Utag1/Uih  ( .x(\Utag1/nh ), .a(ic_itag[6]) );
    inv_1 \Utag1/Uil  ( .x(\Utag1/nl ), .a(ic_itag[1]) );
    ao23_1 \Utag1/Ucl/U1/U1  ( .x(ic_itag[1]), .a(n11), .b(ic_itag[1]), .c(n9), 
        .d(\Utag1/ni ), .e(\Utag1/nh ) );
    ao23_1 \Utag1/Uch/U1/U1  ( .x(ic_itag[6]), .a(n11), .b(ic_itag[6]), .c(n9), 
        .d(tag_id[1]), .e(\Utag1/nl ) );
    inv_1 \Utag0/Uii  ( .x(\Utag0/ni ), .a(tag_id[0]) );
    inv_1 \Utag0/Uih  ( .x(\Utag0/nh ), .a(ic_itag[5]) );
    inv_1 \Utag0/Uil  ( .x(\Utag0/nl ), .a(ic_itag[0]) );
    ao23_1 \Utag0/Ucl/U1/U1  ( .x(ic_itag[0]), .a(n11), .b(ic_itag[0]), .c(n8), 
        .d(\Utag0/ni ), .e(\Utag0/nh ) );
    ao23_1 \Utag0/Uch/U1/U1  ( .x(ic_itag[5]), .a(n10), .b(ic_itag[5]), .c(n8), 
        .d(tag_id[0]), .e(\Utag0/nl ) );
    inv_1 \Usze1/Uii  ( .x(\Usze1/ni ), .a(\size[1] ) );
    inv_1 \Usze1/Uih  ( .x(\Usze1/nh ), .a(ic_size[3]) );
    inv_1 \Usze1/Uil  ( .x(\Usze1/nl ), .a(ic_size[1]) );
    ao23_1 \Usze1/Ucl/U1/U1  ( .x(ic_size[1]), .a(n10), .b(ic_size[1]), .c(n9), 
        .d(\Usze1/ni ), .e(\Usze1/nh ) );
    ao23_1 \Usze1/Uch/U1/U1  ( .x(ic_size[3]), .a(n10), .b(ic_size[3]), .c(n9), 
        .d(\size[1] ), .e(\Usze1/nl ) );
    inv_1 \Usze0/Uii  ( .x(\Usze0/ni ), .a(\size[0] ) );
    inv_1 \Usze0/Uih  ( .x(\Usze0/nh ), .a(ic_size[2]) );
    inv_1 \Usze0/Uil  ( .x(\Usze0/nl ), .a(ic_size[0]) );
    ao23_1 \Usze0/Ucl/U1/U1  ( .x(ic_size[0]), .a(n10), .b(ic_size[0]), .c(n9), 
        .d(\Usze0/ni ), .e(\Usze0/nh ) );
    ao23_1 \Usze0/Uch/U1/U1  ( .x(ic_size[2]), .a(n10), .b(ic_size[2]), .c(n9), 
        .d(\size[0] ), .e(\Usze0/nl ) );
    inv_1 \Urnw/Uii  ( .x(\Urnw/ni ), .a(_24_net_) );
    inv_1 \Urnw/Uih  ( .x(\Urnw/nh ), .a(ic_rnw[1]) );
    inv_1 \Urnw/Uil  ( .x(\Urnw/nl ), .a(ic_rnw[0]) );
    ao23_1 \Urnw/Ucl/U1/U1  ( .x(ic_rnw[0]), .a(n10), .b(ic_rnw[0]), .c(n9), 
        .d(\Urnw/ni ), .e(\Urnw/nh ) );
    ao23_1 \Urnw/Uch/U1/U1  ( .x(ic_rnw[1]), .a(n10), .b(ic_rnw[1]), .c(n9), 
        .d(_24_net_), .e(\Urnw/nl ) );
    inv_1 \Ulock/Uii  ( .x(\Ulock/ni ), .a(mult_o) );
    inv_1 \Ulock/Uih  ( .x(\Ulock/nh ), .a(ic_lock[1]) );
    inv_1 \Ulock/Uil  ( .x(\Ulock/nl ), .a(ic_lock[0]) );
    ao23_1 \Ulock/Ucl/U1/U1  ( .x(ic_lock[0]), .a(n11), .b(ic_lock[0]), .c(n9), 
        .d(\Ulock/ni ), .e(\Ulock/nh ) );
    ao23_1 \Ulock/Uch/U1/U1  ( .x(ic_lock[1]), .a(n11), .b(ic_lock[1]), .c(n8), 
        .d(mult_o), .e(\Ulock/nl ) );
    inv_1 \Upred/Uii  ( .x(\Upred/ni ), .a(prd_o) );
    inv_1 \Upred/Uih  ( .x(\Upred/nh ), .a(ic_pred[1]) );
    inv_1 \Upred/Uil  ( .x(\Upred/nl ), .a(ic_pred[0]) );
    ao23_1 \Upred/Ucl/U1/U1  ( .x(ic_pred[0]), .a(n11), .b(ic_pred[0]), .c(n8), 
        .d(\Upred/ni ), .e(\Upred/nh ) );
    ao23_1 \Upred/Uch/U1/U1  ( .x(ic_pred[1]), .a(n10), .b(ic_pred[1]), .c(n8), 
        .d(prd_o), .e(\Upred/nl ) );
    inv_1 \Useq/Uii  ( .x(\Useq/ni ), .a(seq_o) );
    inv_1 \Useq/Uih  ( .x(\Useq/nh ), .a(ic_seq[1]) );
    inv_1 \Useq/Uil  ( .x(\Useq/nl ), .a(ic_seq[0]) );
    ao23_1 \Useq/Ucl/U1/U1  ( .x(ic_seq[0]), .a(n10), .b(ic_seq[0]), .c(n8), 
        .d(\Useq/ni ), .e(\Useq/nh ) );
    ao23_1 \Useq/Uch/U1/U1  ( .x(ic_seq[1]), .a(n11), .b(ic_seq[1]), .c(n8), 
        .d(seq_o), .e(\Useq/nl ) );
    buf_3 U1 ( .x(n1), .a(en) );
    buf_3 U47 ( .x(n7), .a(en) );
    buf_3 U59 ( .x(n6), .a(en) );
    inv_2 U102 ( .x(n214), .a(n308) );
    inv_0 U112 ( .x(n78), .a(ir_err[0]) );
    nand2i_0 U279 ( .x(_28_net_), .a(ir_err[1]), .b(n72) );
    nand2i_0 U280 ( .x(_25_net_), .a(ir_err[1]), .b(n78) );
    buf_16 U281 ( .x(n8), .a(req_in_delayed) );
    buf_16 U282 ( .x(n9), .a(req_in_delayed) );
    buf_16 U283 ( .x(n10), .a(req_in_delayed) );
    buf_16 U284 ( .x(n11), .a(req_in_delayed) );
endmodule


module master_if_tic ( nReset, mc_req, mc_we, mc_mult, mc_prd, mc_seq, mc_ts, 
    mc_sel, mc_adr, mc_dat, mc_ack, mr_req, mr_we, mr_err, mr_rty, mr_acc, 
    mr_ts, mr_sel, mr_dat, mr_ack, chaincommand, nchaincommandack, 
    chainresponse, nchainresponseack, e_bare, e_dm, e_im, e_wish, r_bare, r_dm, 
    r_im, r_wish, tag_id, force_bare );
input  [2:0] mc_ts;
input  [3:0] mc_sel;
input  [31:0] mc_adr;
input  [31:0] mc_dat;
output [2:0] mr_ts;
output [3:0] mr_sel;
output [31:0] mr_dat;
output [4:0] chaincommand;
input  [4:0] chainresponse;
input  [3:0] e_bare;
input  [3:0] e_dm;
input  [3:0] e_im;
input  [3:0] e_wish;
input  [3:0] r_bare;
input  [3:0] r_dm;
input  [3:0] r_im;
input  [3:0] r_wish;
input  [4:0] tag_id;
input  nReset, mc_req, mc_we, mc_mult, mc_prd, mc_seq, mr_ack, 
    nchaincommandack, force_bare;
output mc_ack, mr_req, mr_we, mr_err, mr_rty, mr_acc, nchainresponseack;
    wire \ci_seq[1] , \ci_seq[0] , \ci_lock[1] , \ci_lock[0] , \ci_rnw[1] , 
        \ci_rnw[0] , \ci_size[3] , \ci_size[2] , \ci_size[1] , \ci_size[0] , 
        \ci_itag[9] , \ci_itag[8] , \ci_itag[7] , \ci_itag[6] , \ci_itag[5] , 
        \ci_itag[4] , \ci_itag[3] , \ci_itag[2] , \ci_itag[1] , \ci_itag[0] , 
        \ci_a[63] , \ci_a[62] , \ci_a[61] , \ci_a[60] , \ci_a[59] , \ci_a[58] , 
        \ci_a[57] , \ci_a[56] , \ci_a[55] , \ci_a[54] , \ci_a[53] , \ci_a[52] , 
        \ci_a[51] , \ci_a[50] , \ci_a[49] , \ci_a[48] , \ci_a[47] , \ci_a[46] , 
        \ci_a[45] , \ci_a[44] , \ci_a[43] , \ci_a[42] , \ci_a[41] , \ci_a[40] , 
        \ci_a[39] , \ci_a[38] , \ci_a[37] , \ci_a[36] , \ci_a[35] , \ci_a[34] , 
        \ci_a[33] , \ci_a[32] , \ci_a[31] , \ci_a[30] , \ci_a[29] , \ci_a[28] , 
        \ci_a[27] , \ci_a[26] , \ci_a[25] , \ci_a[24] , \ci_a[23] , \ci_a[22] , 
        \ci_a[21] , \ci_a[20] , \ci_a[19] , \ci_a[18] , \ci_a[17] , \ci_a[16] , 
        \ci_a[15] , \ci_a[14] , \ci_a[13] , \ci_a[12] , \ci_a[11] , \ci_a[10] , 
        \ci_a[9] , \ci_a[8] , \ci_a[7] , \ci_a[6] , \ci_a[5] , \ci_a[4] , 
        \ci_a[3] , \ci_a[2] , \ci_a[1] , \ci_a[0] , \ci_wd[63] , \ci_wd[62] , 
        \ci_wd[61] , \ci_wd[60] , \ci_wd[59] , \ci_wd[58] , \ci_wd[57] , 
        \ci_wd[56] , \ci_wd[55] , \ci_wd[54] , \ci_wd[53] , \ci_wd[52] , 
        \ci_wd[51] , \ci_wd[50] , \ci_wd[49] , \ci_wd[48] , \ci_wd[47] , 
        \ci_wd[46] , \ci_wd[45] , \ci_wd[44] , \ci_wd[43] , \ci_wd[42] , 
        \ci_wd[41] , \ci_wd[40] , \ci_wd[39] , \ci_wd[38] , \ci_wd[37] , 
        \ci_wd[36] , \ci_wd[35] , \ci_wd[34] , \ci_wd[33] , \ci_wd[32] , 
        \ci_wd[31] , \ci_wd[30] , \ci_wd[29] , \ci_wd[28] , \ci_wd[27] , 
        \ci_wd[26] , \ci_wd[25] , \ci_wd[24] , \ci_wd[23] , \ci_wd[22] , 
        \ci_wd[21] , \ci_wd[20] , \ci_wd[19] , \ci_wd[18] , \ci_wd[17] , 
        \ci_wd[16] , \ci_wd[15] , \ci_wd[14] , \ci_wd[13] , \ci_wd[12] , 
        \ci_wd[11] , \ci_wd[10] , \ci_wd[9] , \ci_wd[8] , \ci_wd[7] , 
        \ci_wd[6] , \ci_wd[5] , \ci_wd[4] , \ci_wd[3] , \ci_wd[2] , \ci_wd[1] , 
        \ci_wd[0] , \ci_pred[1] , \ci_pred[0] , \ci_col[5] , \ci_col[4] , 
        \ci_col[3] , \ci_col[2] , \ci_col[1] , \ci_col[0] , ci_ack, 
        \ri_err[1] , \ri_err[0] , \ri_rnw[1] , \ri_rnw[0] , \ri_rd[63] , 
        \ri_rd[62] , \ri_rd[61] , \ri_rd[60] , \ri_rd[59] , \ri_rd[58] , 
        \ri_rd[57] , \ri_rd[56] , \ri_rd[55] , \ri_rd[54] , \ri_rd[53] , 
        \ri_rd[52] , \ri_rd[51] , \ri_rd[50] , \ri_rd[49] , \ri_rd[48] , 
        \ri_rd[47] , \ri_rd[46] , \ri_rd[45] , \ri_rd[44] , \ri_rd[43] , 
        \ri_rd[42] , \ri_rd[41] , \ri_rd[40] , \ri_rd[39] , \ri_rd[38] , 
        \ri_rd[37] , \ri_rd[36] , \ri_rd[35] , \ri_rd[34] , \ri_rd[33] , 
        \ri_rd[32] , \ri_rd[31] , \ri_rd[30] , \ri_rd[29] , \ri_rd[28] , 
        \ri_rd[27] , \ri_rd[26] , \ri_rd[25] , \ri_rd[24] , \ri_rd[23] , 
        \ri_rd[22] , \ri_rd[21] , \ri_rd[20] , \ri_rd[19] , \ri_rd[18] , 
        \ri_rd[17] , \ri_rd[16] , \ri_rd[15] , \ri_rd[14] , \ri_rd[13] , 
        \ri_rd[12] , \ri_rd[11] , \ri_rd[10] , \ri_rd[9] , \ri_rd[8] , 
        \ri_rd[7] , \ri_rd[6] , \ri_rd[5] , \ri_rd[4] , \ri_rd[3] , \ri_rd[2] , 
        \ri_rd[1] , \ri_rd[0] , ri_ack, reset, nroute_ack, routetx_req, 
        routetx_ack, \route[4] , \route[1] , \route[0] , \i_eh[2] , \i_eh[1] , 
        \i_eh[0] , \i_el[3] , \i_el[2] , \i_el[1] , \i_el[0] , \i_rh[3] , 
        \i_rh[2] , \i_rh[1] , \i_rl[3] , \i_rl[2] , \i_rl[1] , \i_rl[0] ;
    wire SYNOPSYS_UNCONNECTED_1 , SYNOPSYS_UNCONNECTED_2 , 
	SYNOPSYS_UNCONNECTED_3 , SYNOPSYS_UNCONNECTED_4 ;
    assign mr_rty = 1'b0;
    assign mr_acc = 1'b0;
    assign mr_ts[2] = 1'b0;
    assign mr_ts[1] = 1'b0;
    assign mr_ts[0] = 1'b0;
    inv_2 U1 ( .x(reset), .a(nReset) );
    m2cp_tic master2chainif ( .req_in(mc_req), .ts_o(mc_ts), .sel_o(mc_sel), 
        .mult_o(mc_mult), .we_o(mc_we), .prd_o(mc_prd), .seq_o(mc_seq), 
        .adr_o(mc_adr), .dat_o(mc_dat), .ain(mc_ack), .ic_seq({\ci_seq[1] , 
        \ci_seq[0] }), .ic_pred({\ci_pred[1] , \ci_pred[0] }), .ic_size({
        \ci_size[3] , \ci_size[2] , \ci_size[1] , \ci_size[0] }), .ic_itag({
        \ci_itag[9] , \ci_itag[8] , \ci_itag[7] , \ci_itag[6] , \ci_itag[5] , 
        \ci_itag[4] , \ci_itag[3] , \ci_itag[2] , \ci_itag[1] , \ci_itag[0] }), 
        .ic_wd({\ci_wd[63] , \ci_wd[62] , \ci_wd[61] , \ci_wd[60] , 
        \ci_wd[59] , \ci_wd[58] , \ci_wd[57] , \ci_wd[56] , \ci_wd[55] , 
        \ci_wd[54] , \ci_wd[53] , \ci_wd[52] , \ci_wd[51] , \ci_wd[50] , 
        \ci_wd[49] , \ci_wd[48] , \ci_wd[47] , \ci_wd[46] , \ci_wd[45] , 
        \ci_wd[44] , \ci_wd[43] , \ci_wd[42] , \ci_wd[41] , \ci_wd[40] , 
        \ci_wd[39] , \ci_wd[38] , \ci_wd[37] , \ci_wd[36] , \ci_wd[35] , 
        \ci_wd[34] , \ci_wd[33] , \ci_wd[32] , \ci_wd[31] , \ci_wd[30] , 
        \ci_wd[29] , \ci_wd[28] , \ci_wd[27] , \ci_wd[26] , \ci_wd[25] , 
        \ci_wd[24] , \ci_wd[23] , \ci_wd[22] , \ci_wd[21] , \ci_wd[20] , 
        \ci_wd[19] , \ci_wd[18] , \ci_wd[17] , \ci_wd[16] , \ci_wd[15] , 
        \ci_wd[14] , \ci_wd[13] , \ci_wd[12] , \ci_wd[11] , \ci_wd[10] , 
        \ci_wd[9] , \ci_wd[8] , \ci_wd[7] , \ci_wd[6] , \ci_wd[5] , \ci_wd[4] , 
        \ci_wd[3] , \ci_wd[2] , \ci_wd[1] , \ci_wd[0] }), .ic_lock({
        \ci_lock[1] , \ci_lock[0] }), .ic_a({\ci_a[63] , \ci_a[62] , 
        \ci_a[61] , \ci_a[60] , \ci_a[59] , \ci_a[58] , \ci_a[57] , \ci_a[56] , 
        \ci_a[55] , \ci_a[54] , \ci_a[53] , \ci_a[52] , \ci_a[51] , \ci_a[50] , 
        \ci_a[49] , \ci_a[48] , \ci_a[47] , \ci_a[46] , \ci_a[45] , \ci_a[44] , 
        \ci_a[43] , \ci_a[42] , \ci_a[41] , \ci_a[40] , \ci_a[39] , \ci_a[38] , 
        \ci_a[37] , \ci_a[36] , \ci_a[35] , \ci_a[34] , \ci_a[33] , \ci_a[32] , 
        \ci_a[31] , \ci_a[30] , \ci_a[29] , \ci_a[28] , \ci_a[27] , \ci_a[26] , 
        \ci_a[25] , \ci_a[24] , \ci_a[23] , \ci_a[22] , \ci_a[21] , \ci_a[20] , 
        \ci_a[19] , \ci_a[18] , \ci_a[17] , \ci_a[16] , \ci_a[15] , \ci_a[14] , 
        \ci_a[13] , \ci_a[12] , \ci_a[11] , \ci_a[10] , \ci_a[9] , \ci_a[8] , 
        \ci_a[7] , \ci_a[6] , \ci_a[5] , \ci_a[4] , \ci_a[3] , \ci_a[2] , 
        \ci_a[1] , \ci_a[0] }), .ic_rnw({\ci_rnw[1] , \ci_rnw[0] }), .ic_col({
        \ci_col[5] , \ci_col[4] , \ci_col[3] , \ci_col[2] , \ci_col[1] , 
        \ci_col[0] }), .ic_ack(ci_ack), .req_out(mr_req), .we_i(mr_we), 
        .err_i(mr_err), .dat_i(mr_dat), .aout(mr_ack), .ir_rd({\ri_rd[63] , 
        \ri_rd[62] , \ri_rd[61] , \ri_rd[60] , \ri_rd[59] , \ri_rd[58] , 
        \ri_rd[57] , \ri_rd[56] , \ri_rd[55] , \ri_rd[54] , \ri_rd[53] , 
        \ri_rd[52] , \ri_rd[51] , \ri_rd[50] , \ri_rd[49] , \ri_rd[48] , 
        \ri_rd[47] , \ri_rd[46] , \ri_rd[45] , \ri_rd[44] , \ri_rd[43] , 
        \ri_rd[42] , \ri_rd[41] , \ri_rd[40] , \ri_rd[39] , \ri_rd[38] , 
        \ri_rd[37] , \ri_rd[36] , \ri_rd[35] , \ri_rd[34] , \ri_rd[33] , 
        \ri_rd[32] , \ri_rd[31] , \ri_rd[30] , \ri_rd[29] , \ri_rd[28] , 
        \ri_rd[27] , \ri_rd[26] , \ri_rd[25] , \ri_rd[24] , \ri_rd[23] , 
        \ri_rd[22] , \ri_rd[21] , \ri_rd[20] , \ri_rd[19] , \ri_rd[18] , 
        \ri_rd[17] , \ri_rd[16] , \ri_rd[15] , \ri_rd[14] , \ri_rd[13] , 
        \ri_rd[12] , \ri_rd[11] , \ri_rd[10] , \ri_rd[9] , \ri_rd[8] , 
        \ri_rd[7] , \ri_rd[6] , \ri_rd[5] , \ri_rd[4] , \ri_rd[3] , \ri_rd[2] , 
        \ri_rd[1] , \ri_rd[0] }), .ir_err({\ri_err[1] , \ri_err[0] }), 
        .ir_rnw({\ri_rnw[1] , \ri_rnw[0] }), .ir_ack(ri_ack), .tag_id(tag_id), 
        .reset(reset) );
    i_adec_tic dec ( .e_h({SYNOPSYS_UNCONNECTED_1, \i_eh[2] , \i_eh[1] , 
        \i_eh[0] }), .e_l({\i_el[3] , \i_el[2] , \i_el[1] , \i_el[0] }), .r_h(
        {\i_rh[3] , \i_rh[2] , \i_rh[1] , SYNOPSYS_UNCONNECTED_2}), .r_l({
        \i_rl[3] , \i_rl[2] , \i_rl[1] , \i_rl[0] }), .ah({\ci_a[63] , 
        \ci_a[62] , \ci_a[61] , \ci_a[60] , \ci_a[59] , \ci_a[58] , \ci_a[57] , 
        \ci_a[56] , \ci_a[55] , \ci_a[54] , \ci_a[53] , \ci_a[52] , \ci_a[51] , 
        \ci_a[50] , \ci_a[49] , \ci_a[48] , \ci_a[47] , \ci_a[46] , \ci_a[45] , 
        \ci_a[44] , \ci_a[43] , \ci_a[42] , \ci_a[41] , \ci_a[40] , \ci_a[39] , 
        \ci_a[38] , \ci_a[37] , \ci_a[36] , \ci_a[35] , \ci_a[34] , \ci_a[33] , 
        \ci_a[32] }), .al({\ci_a[31] , \ci_a[30] , \ci_a[29] , \ci_a[28] , 
        \ci_a[27] , \ci_a[26] , \ci_a[25] , \ci_a[24] , \ci_a[23] , \ci_a[22] , 
        \ci_a[21] , \ci_a[20] , \ci_a[19] , \ci_a[18] , \ci_a[17] , \ci_a[16] , 
        \ci_a[15] , \ci_a[14] , \ci_a[13] , \ci_a[12] , \ci_a[11] , \ci_a[10] , 
        \ci_a[9] , \ci_a[8] , \ci_a[7] , \ci_a[6] , \ci_a[5] , \ci_a[4] , 
        \ci_a[3] , \ci_a[2] , \ci_a[1] , \ci_a[0] }), .e_bare(e_bare), .e_dm(
        e_dm), .e_im(e_im), .e_wish(e_wish), .r_bare(r_bare), .r_dm(r_dm), 
        .r_im(r_im), .r_wish(r_wish), .force_bare(force_bare) );
    route_tx_tic rt ( .o({\route[4] , SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, \route[1] , \route[0] }), .rtxack(routetx_ack), 
        .e_h({1'b0, \i_eh[2] , \i_eh[1] , \i_eh[0] }), .e_l({\i_el[3] , 
        \i_el[2] , \i_el[1] , \i_el[0] }), .noa(nroute_ack), .r_h({\i_rh[3] , 
        \i_rh[2] , \i_rh[1] , 1'b0}), .r_l({\i_rl[3] , \i_rl[2] , \i_rl[1] , 
        \i_rl[0] }), .rtxreq(routetx_req) );
    initiator_tic it ( .cack(ci_ack), .chaincommand(chaincommand), .err({
        \ri_err[1] , \ri_err[0] }), .nchainresponseack(nchainresponseack), 
        .nrouteack(nroute_ack), .rd({\ri_rd[63] , \ri_rd[62] , \ri_rd[61] , 
        \ri_rd[60] , \ri_rd[59] , \ri_rd[58] , \ri_rd[57] , \ri_rd[56] , 
        \ri_rd[55] , \ri_rd[54] , \ri_rd[53] , \ri_rd[52] , \ri_rd[51] , 
        \ri_rd[50] , \ri_rd[49] , \ri_rd[48] , \ri_rd[47] , \ri_rd[46] , 
        \ri_rd[45] , \ri_rd[44] , \ri_rd[43] , \ri_rd[42] , \ri_rd[41] , 
        \ri_rd[40] , \ri_rd[39] , \ri_rd[38] , \ri_rd[37] , \ri_rd[36] , 
        \ri_rd[35] , \ri_rd[34] , \ri_rd[33] , \ri_rd[32] , \ri_rd[31] , 
        \ri_rd[30] , \ri_rd[29] , \ri_rd[28] , \ri_rd[27] , \ri_rd[26] , 
        \ri_rd[25] , \ri_rd[24] , \ri_rd[23] , \ri_rd[22] , \ri_rd[21] , 
        \ri_rd[20] , \ri_rd[19] , \ri_rd[18] , \ri_rd[17] , \ri_rd[16] , 
        \ri_rd[15] , \ri_rd[14] , \ri_rd[13] , \ri_rd[12] , \ri_rd[11] , 
        \ri_rd[10] , \ri_rd[9] , \ri_rd[8] , \ri_rd[7] , \ri_rd[6] , 
        \ri_rd[5] , \ri_rd[4] , \ri_rd[3] , \ri_rd[2] , \ri_rd[1] , \ri_rd[0] 
        }), .routetxreq(routetx_req), .rrnw({\ri_rnw[1] , \ri_rnw[0] }), .a({
        \ci_a[63] , \ci_a[62] , \ci_a[61] , \ci_a[60] , \ci_a[59] , \ci_a[58] , 
        \ci_a[57] , \ci_a[56] , \ci_a[55] , \ci_a[54] , \ci_a[53] , \ci_a[52] , 
        \ci_a[51] , \ci_a[50] , \ci_a[49] , \ci_a[48] , \ci_a[47] , \ci_a[46] , 
        \ci_a[45] , \ci_a[44] , \ci_a[43] , \ci_a[42] , \ci_a[41] , \ci_a[40] , 
        \ci_a[39] , \ci_a[38] , \ci_a[37] , \ci_a[36] , \ci_a[35] , \ci_a[34] , 
        \ci_a[33] , \ci_a[32] , \ci_a[31] , \ci_a[30] , \ci_a[29] , \ci_a[28] , 
        \ci_a[27] , \ci_a[26] , \ci_a[25] , \ci_a[24] , \ci_a[23] , \ci_a[22] , 
        \ci_a[21] , \ci_a[20] , \ci_a[19] , \ci_a[18] , \ci_a[17] , \ci_a[16] , 
        \ci_a[15] , \ci_a[14] , \ci_a[13] , \ci_a[12] , \ci_a[11] , \ci_a[10] , 
        \ci_a[9] , \ci_a[8] , \ci_a[7] , \ci_a[6] , \ci_a[5] , \ci_a[4] , 
        \ci_a[3] , \ci_a[2] , \ci_a[1] , \ci_a[0] }), .chainresponse(
        chainresponse), .col({\ci_col[5] , \ci_col[4] , \ci_col[3] , 
        \ci_col[2] , \ci_col[1] , \ci_col[0] }), .crnw({\ci_rnw[1] , 
        \ci_rnw[0] }), .itag({\ci_itag[9] , \ci_itag[8] , \ci_itag[7] , 
        \ci_itag[6] , \ci_itag[5] , \ci_itag[4] , \ci_itag[3] , \ci_itag[2] , 
        \ci_itag[1] , \ci_itag[0] }), .lock({\ci_lock[1] , \ci_lock[0] }), 
        .nReset(nReset), .nchaincommandack(nchaincommandack), .pred({
        \ci_pred[1] , \ci_pred[0] }), .rack(ri_ack), .route({\route[4] , 1'b0, 
        1'b0, \route[1] , \route[0] }), .routetxack(routetx_ack), .seq({
        \ci_seq[1] , \ci_seq[0] }), .size({\ci_size[3] , \ci_size[2] , 
        \ci_size[1] , \ci_size[0] }), .wd({\ci_wd[63] , \ci_wd[62] , 
        \ci_wd[61] , \ci_wd[60] , \ci_wd[59] , \ci_wd[58] , \ci_wd[57] , 
        \ci_wd[56] , \ci_wd[55] , \ci_wd[54] , \ci_wd[53] , \ci_wd[52] , 
        \ci_wd[51] , \ci_wd[50] , \ci_wd[49] , \ci_wd[48] , \ci_wd[47] , 
        \ci_wd[46] , \ci_wd[45] , \ci_wd[44] , \ci_wd[43] , \ci_wd[42] , 
        \ci_wd[41] , \ci_wd[40] , \ci_wd[39] , \ci_wd[38] , \ci_wd[37] , 
        \ci_wd[36] , \ci_wd[35] , \ci_wd[34] , \ci_wd[33] , \ci_wd[32] , 
        \ci_wd[31] , \ci_wd[30] , \ci_wd[29] , \ci_wd[28] , \ci_wd[27] , 
        \ci_wd[26] , \ci_wd[25] , \ci_wd[24] , \ci_wd[23] , \ci_wd[22] , 
        \ci_wd[21] , \ci_wd[20] , \ci_wd[19] , \ci_wd[18] , \ci_wd[17] , 
        \ci_wd[16] , \ci_wd[15] , \ci_wd[14] , \ci_wd[13] , \ci_wd[12] , 
        \ci_wd[11] , \ci_wd[10] , \ci_wd[9] , \ci_wd[8] , \ci_wd[7] , 
        \ci_wd[6] , \ci_wd[5] , \ci_wd[4] , \ci_wd[3] , \ci_wd[2] , \ci_wd[1] , 
        \ci_wd[0] }) );
endmodule


module t_adec_imem ( e_h, e_l, r_h, r_l, e_dp, e_ip, e_tic, r_dp, r_ip, r_tic, 
    tag_h, tag_l );
output [2:0] e_h;
output [2:0] e_l;
output [2:0] r_h;
output [2:0] r_l;
input  [2:0] e_dp;
input  [2:0] e_ip;
input  [2:0] e_tic;
input  [2:0] r_dp;
input  [2:0] r_ip;
input  [2:0] r_tic;
input  [4:0] tag_h;
input  [4:0] tag_l;
    wire \e_l[2] , \e_l[1] , \tag_h[4] , \e_l[0] ;
    assign e_h[2] = 1'b0;
    assign e_h[1] = \e_l[0] ;
    assign e_h[0] = \e_l[1] ;
    assign e_l[2] = \e_l[2] ;
    assign e_l[1] = \e_l[1] ;
    assign e_l[0] = \e_l[0] ;
    assign r_h[2] = \e_l[1] ;
    assign r_h[1] = \tag_h[4] ;
    assign r_h[0] = 1'b0;
    assign r_l[2] = \e_l[0] ;
    assign r_l[0] = \e_l[2] ;
    assign \tag_h[4]  = tag_h[4];
    or2_1 U3 ( .x(r_l[1]), .a(\e_l[0] ), .b(tag_h[3]) );
    buf_3 U6 ( .x(\e_l[0] ), .a(tag_h[2]) );
    or2_2 U7 ( .x(\e_l[2] ), .a(\tag_h[4] ), .b(r_l[1]) );
    or2_2 U8 ( .x(\e_l[1] ), .a(tag_h[3]), .b(\tag_h[4] ) );
endmodule


module chain_sendmux8_8 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/naa , \U1693/bdone , \U1693/net3 , 
        \U1693/drivemonitor , \U1693/net2 , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendmux8_9 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/naa , \U1693/bdone , \U1693/net3 , 
        \U1693/drivemonitor , \U1693/net2 , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendmux8_10 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/naa , \U1693/bdone , \U1693/net3 , 
        \U1693/drivemonitor , \U1693/net2 , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendmux8_11 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/naa , \U1693/bdone , \U1693/net3 , 
        \U1693/drivemonitor , \U1693/net2 , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendword_1 ( ctrlack, oh, ol, chainackff, ctrlreq, ih, il );
output [7:0] oh;
output [7:0] ol;
input  [31:0] ih;
input  [31:0] il;
input  chainackff, ctrlreq;
output ctrlack;
    wire \third_oh[7] , \third_oh[6] , \third_oh[5] , \third_oh[4] , 
        \third_oh[3] , \third_oh[2] , \third_oh[1] , \third_oh[0] , 
        \fourth_ol[7] , \fourth_ol[6] , \fourth_ol[5] , \fourth_ol[4] , 
        \fourth_ol[3] , \fourth_ol[2] , \fourth_ol[1] , \fourth_ol[0] , 
        \third_ol[7] , \third_ol[6] , \third_ol[5] , \third_ol[4] , 
        \third_ol[3] , \third_ol[2] , \third_ol[1] , \third_ol[0] , 
        \fourth_oh[7] , \fourth_oh[6] , \fourth_oh[5] , \fourth_oh[4] , 
        \fourth_oh[3] , \fourth_oh[2] , \fourth_oh[1] , \fourth_oh[0] , 
        \second_oh[7] , \second_oh[6] , \second_oh[5] , \second_oh[4] , 
        \second_oh[3] , \second_oh[2] , \second_oh[1] , \second_oh[0] , 
        \second_ol[7] , \second_ol[6] , \second_ol[5] , \second_ol[4] , 
        \second_ol[3] , \second_ol[2] , \second_ol[1] , \second_ol[0] , 
        \first_oh[7] , \first_oh[6] , \first_oh[5] , \first_oh[4] , 
        \first_oh[3] , \first_oh[2] , \first_oh[1] , \first_oh[0] , 
        \first_ol[7] , \first_ol[6] , \first_ol[5] , \first_ol[4] , 
        \first_ol[3] , \first_ol[2] , \first_ol[1] , \first_ol[0] , net44, 
        net51, net58, bctrlreq, \U309_0_/n5 , \U309_0_/n1 , \U309_0_/n2 , 
        \U309_0_/n3 , \U309_0_/n4 , \U309_1_/n5 , \U309_1_/n1 , \U309_1_/n2 , 
        \U309_1_/n3 , \U309_1_/n4 , \U309_2_/n5 , \U309_2_/n1 , \U309_2_/n2 , 
        \U309_2_/n3 , \U309_2_/n4 , \U309_3_/n5 , \U309_3_/n1 , \U309_3_/n2 , 
        \U309_3_/n3 , \U309_3_/n4 , \U309_4_/n5 , \U309_4_/n1 , \U309_4_/n2 , 
        \U309_4_/n3 , \U309_4_/n4 , \U309_5_/n5 , \U309_5_/n1 , \U309_5_/n2 , 
        \U309_5_/n3 , \U309_5_/n4 , \U309_6_/n5 , \U309_6_/n1 , \U309_6_/n2 , 
        \U309_6_/n3 , \U309_6_/n4 , \U309_7_/n5 , \U309_7_/n1 , \U309_7_/n2 , 
        \U309_7_/n3 , \U309_7_/n4 , \U310_0_/n5 , \U310_0_/n1 , \U310_0_/n2 , 
        \U310_0_/n3 , \U310_0_/n4 , \U310_1_/n5 , \U310_1_/n1 , \U310_1_/n2 , 
        \U310_1_/n3 , \U310_1_/n4 , \U310_2_/n5 , \U310_2_/n1 , \U310_2_/n2 , 
        \U310_2_/n3 , \U310_2_/n4 , \U310_3_/n5 , \U310_3_/n1 , \U310_3_/n2 , 
        \U310_3_/n3 , \U310_3_/n4 , \U310_4_/n5 , \U310_4_/n1 , \U310_4_/n2 , 
        \U310_4_/n3 , \U310_4_/n4 , \U310_5_/n5 , \U310_5_/n1 , \U310_5_/n2 , 
        \U310_5_/n3 , \U310_5_/n4 , \U310_6_/n5 , \U310_6_/n1 , \U310_6_/n2 , 
        \U310_6_/n3 , \U310_6_/n4 , \U310_7_/n5 , \U310_7_/n1 , \U310_7_/n2 , 
        \U310_7_/n3 , \U310_7_/n4 ;
    chain_sendmux8_10 I4 ( .ctrlack(ctrlack), .oh({\fourth_oh[7] , 
        \fourth_oh[6] , \fourth_oh[5] , \fourth_oh[4] , \fourth_oh[3] , 
        \fourth_oh[2] , \fourth_oh[1] , \fourth_oh[0] }), .ol({\fourth_ol[7] , 
        \fourth_ol[6] , \fourth_ol[5] , \fourth_ol[4] , \fourth_ol[3] , 
        \fourth_ol[2] , \fourth_ol[1] , \fourth_ol[0] }), .i_h(ih[7:0]), .i_l(
        il[7:0]), .ctrlreq(net44), .oa(chainackff) );
    chain_sendmux8_9 I3 ( .ctrlack(net44), .oh({\third_oh[7] , \third_oh[6] , 
        \third_oh[5] , \third_oh[4] , \third_oh[3] , \third_oh[2] , 
        \third_oh[1] , \third_oh[0] }), .ol({\third_ol[7] , \third_ol[6] , 
        \third_ol[5] , \third_ol[4] , \third_ol[3] , \third_ol[2] , 
        \third_ol[1] , \third_ol[0] }), .i_h(ih[15:8]), .i_l(il[15:8]), 
        .ctrlreq(net51), .oa(chainackff) );
    chain_sendmux8_8 I2 ( .ctrlack(net51), .oh({\second_oh[7] , \second_oh[6] , 
        \second_oh[5] , \second_oh[4] , \second_oh[3] , \second_oh[2] , 
        \second_oh[1] , \second_oh[0] }), .ol({\second_ol[7] , \second_ol[6] , 
        \second_ol[5] , \second_ol[4] , \second_ol[3] , \second_ol[2] , 
        \second_ol[1] , \second_ol[0] }), .i_h(ih[23:16]), .i_l(il[23:16]), 
        .ctrlreq(net58), .oa(chainackff) );
    chain_sendmux8_11 U320 ( .ctrlack(net58), .oh({\first_oh[7] , 
        \first_oh[6] , \first_oh[5] , \first_oh[4] , \first_oh[3] , 
        \first_oh[2] , \first_oh[1] , \first_oh[0] }), .ol({\first_ol[7] , 
        \first_ol[6] , \first_ol[5] , \first_ol[4] , \first_ol[3] , 
        \first_ol[2] , \first_ol[1] , \first_ol[0] }), .i_h(ih[31:24]), .i_l(
        il[31:24]), .ctrlreq(bctrlreq), .oa(chainackff) );
    buf_2 \U328/U7  ( .x(bctrlreq), .a(ctrlreq) );
    and4_2 \U309_0_/U24  ( .x(\U309_0_/n5 ), .a(\U309_0_/n1 ), .b(\U309_0_/n2 
        ), .c(\U309_0_/n3 ), .d(\U309_0_/n4 ) );
    inv_1 \U309_0_/U1  ( .x(\U309_0_/n1 ), .a(\fourth_oh[0] ) );
    inv_1 \U309_0_/U2  ( .x(\U309_0_/n2 ), .a(\third_oh[0] ) );
    inv_1 \U309_0_/U3  ( .x(\U309_0_/n3 ), .a(\second_oh[0] ) );
    inv_1 \U309_0_/U4  ( .x(\U309_0_/n4 ), .a(\first_oh[0] ) );
    inv_4 \U309_0_/U5  ( .x(oh[0]), .a(\U309_0_/n5 ) );
    and4_2 \U309_1_/U24  ( .x(\U309_1_/n5 ), .a(\U309_1_/n1 ), .b(\U309_1_/n2 
        ), .c(\U309_1_/n3 ), .d(\U309_1_/n4 ) );
    inv_1 \U309_1_/U1  ( .x(\U309_1_/n1 ), .a(\fourth_oh[1] ) );
    inv_1 \U309_1_/U2  ( .x(\U309_1_/n2 ), .a(\third_oh[1] ) );
    inv_1 \U309_1_/U3  ( .x(\U309_1_/n3 ), .a(\second_oh[1] ) );
    inv_1 \U309_1_/U4  ( .x(\U309_1_/n4 ), .a(\first_oh[1] ) );
    inv_4 \U309_1_/U5  ( .x(oh[1]), .a(\U309_1_/n5 ) );
    and4_2 \U309_2_/U24  ( .x(\U309_2_/n5 ), .a(\U309_2_/n1 ), .b(\U309_2_/n2 
        ), .c(\U309_2_/n3 ), .d(\U309_2_/n4 ) );
    inv_1 \U309_2_/U1  ( .x(\U309_2_/n1 ), .a(\fourth_oh[2] ) );
    inv_1 \U309_2_/U2  ( .x(\U309_2_/n2 ), .a(\third_oh[2] ) );
    inv_1 \U309_2_/U3  ( .x(\U309_2_/n3 ), .a(\second_oh[2] ) );
    inv_1 \U309_2_/U4  ( .x(\U309_2_/n4 ), .a(\first_oh[2] ) );
    inv_4 \U309_2_/U5  ( .x(oh[2]), .a(\U309_2_/n5 ) );
    and4_2 \U309_3_/U24  ( .x(\U309_3_/n5 ), .a(\U309_3_/n1 ), .b(\U309_3_/n2 
        ), .c(\U309_3_/n3 ), .d(\U309_3_/n4 ) );
    inv_1 \U309_3_/U1  ( .x(\U309_3_/n1 ), .a(\fourth_oh[3] ) );
    inv_1 \U309_3_/U2  ( .x(\U309_3_/n2 ), .a(\third_oh[3] ) );
    inv_1 \U309_3_/U3  ( .x(\U309_3_/n3 ), .a(\second_oh[3] ) );
    inv_1 \U309_3_/U4  ( .x(\U309_3_/n4 ), .a(\first_oh[3] ) );
    inv_4 \U309_3_/U5  ( .x(oh[3]), .a(\U309_3_/n5 ) );
    and4_2 \U309_4_/U24  ( .x(\U309_4_/n5 ), .a(\U309_4_/n1 ), .b(\U309_4_/n2 
        ), .c(\U309_4_/n3 ), .d(\U309_4_/n4 ) );
    inv_1 \U309_4_/U1  ( .x(\U309_4_/n1 ), .a(\fourth_oh[4] ) );
    inv_1 \U309_4_/U2  ( .x(\U309_4_/n2 ), .a(\third_oh[4] ) );
    inv_1 \U309_4_/U3  ( .x(\U309_4_/n3 ), .a(\second_oh[4] ) );
    inv_1 \U309_4_/U4  ( .x(\U309_4_/n4 ), .a(\first_oh[4] ) );
    inv_4 \U309_4_/U5  ( .x(oh[4]), .a(\U309_4_/n5 ) );
    and4_2 \U309_5_/U24  ( .x(\U309_5_/n5 ), .a(\U309_5_/n1 ), .b(\U309_5_/n2 
        ), .c(\U309_5_/n3 ), .d(\U309_5_/n4 ) );
    inv_1 \U309_5_/U1  ( .x(\U309_5_/n1 ), .a(\fourth_oh[5] ) );
    inv_1 \U309_5_/U2  ( .x(\U309_5_/n2 ), .a(\third_oh[5] ) );
    inv_1 \U309_5_/U3  ( .x(\U309_5_/n3 ), .a(\second_oh[5] ) );
    inv_1 \U309_5_/U4  ( .x(\U309_5_/n4 ), .a(\first_oh[5] ) );
    inv_4 \U309_5_/U5  ( .x(oh[5]), .a(\U309_5_/n5 ) );
    and4_2 \U309_6_/U24  ( .x(\U309_6_/n5 ), .a(\U309_6_/n1 ), .b(\U309_6_/n2 
        ), .c(\U309_6_/n3 ), .d(\U309_6_/n4 ) );
    inv_1 \U309_6_/U1  ( .x(\U309_6_/n1 ), .a(\fourth_oh[6] ) );
    inv_1 \U309_6_/U2  ( .x(\U309_6_/n2 ), .a(\third_oh[6] ) );
    inv_1 \U309_6_/U3  ( .x(\U309_6_/n3 ), .a(\second_oh[6] ) );
    inv_1 \U309_6_/U4  ( .x(\U309_6_/n4 ), .a(\first_oh[6] ) );
    inv_4 \U309_6_/U5  ( .x(oh[6]), .a(\U309_6_/n5 ) );
    and4_2 \U309_7_/U24  ( .x(\U309_7_/n5 ), .a(\U309_7_/n1 ), .b(\U309_7_/n2 
        ), .c(\U309_7_/n3 ), .d(\U309_7_/n4 ) );
    inv_1 \U309_7_/U1  ( .x(\U309_7_/n1 ), .a(\fourth_oh[7] ) );
    inv_1 \U309_7_/U2  ( .x(\U309_7_/n2 ), .a(\third_oh[7] ) );
    inv_1 \U309_7_/U3  ( .x(\U309_7_/n3 ), .a(\second_oh[7] ) );
    inv_1 \U309_7_/U4  ( .x(\U309_7_/n4 ), .a(\first_oh[7] ) );
    inv_4 \U309_7_/U5  ( .x(oh[7]), .a(\U309_7_/n5 ) );
    and4_2 \U310_0_/U24  ( .x(\U310_0_/n5 ), .a(\U310_0_/n1 ), .b(\U310_0_/n2 
        ), .c(\U310_0_/n3 ), .d(\U310_0_/n4 ) );
    inv_1 \U310_0_/U1  ( .x(\U310_0_/n1 ), .a(\fourth_ol[0] ) );
    inv_1 \U310_0_/U2  ( .x(\U310_0_/n2 ), .a(\third_ol[0] ) );
    inv_1 \U310_0_/U3  ( .x(\U310_0_/n3 ), .a(\second_ol[0] ) );
    inv_1 \U310_0_/U4  ( .x(\U310_0_/n4 ), .a(\first_ol[0] ) );
    inv_4 \U310_0_/U5  ( .x(ol[0]), .a(\U310_0_/n5 ) );
    and4_2 \U310_1_/U24  ( .x(\U310_1_/n5 ), .a(\U310_1_/n1 ), .b(\U310_1_/n2 
        ), .c(\U310_1_/n3 ), .d(\U310_1_/n4 ) );
    inv_1 \U310_1_/U1  ( .x(\U310_1_/n1 ), .a(\fourth_ol[1] ) );
    inv_1 \U310_1_/U2  ( .x(\U310_1_/n2 ), .a(\third_ol[1] ) );
    inv_1 \U310_1_/U3  ( .x(\U310_1_/n3 ), .a(\second_ol[1] ) );
    inv_1 \U310_1_/U4  ( .x(\U310_1_/n4 ), .a(\first_ol[1] ) );
    inv_4 \U310_1_/U5  ( .x(ol[1]), .a(\U310_1_/n5 ) );
    and4_2 \U310_2_/U24  ( .x(\U310_2_/n5 ), .a(\U310_2_/n1 ), .b(\U310_2_/n2 
        ), .c(\U310_2_/n3 ), .d(\U310_2_/n4 ) );
    inv_1 \U310_2_/U1  ( .x(\U310_2_/n1 ), .a(\fourth_ol[2] ) );
    inv_1 \U310_2_/U2  ( .x(\U310_2_/n2 ), .a(\third_ol[2] ) );
    inv_1 \U310_2_/U3  ( .x(\U310_2_/n3 ), .a(\second_ol[2] ) );
    inv_1 \U310_2_/U4  ( .x(\U310_2_/n4 ), .a(\first_ol[2] ) );
    inv_4 \U310_2_/U5  ( .x(ol[2]), .a(\U310_2_/n5 ) );
    and4_2 \U310_3_/U24  ( .x(\U310_3_/n5 ), .a(\U310_3_/n1 ), .b(\U310_3_/n2 
        ), .c(\U310_3_/n3 ), .d(\U310_3_/n4 ) );
    inv_1 \U310_3_/U1  ( .x(\U310_3_/n1 ), .a(\fourth_ol[3] ) );
    inv_1 \U310_3_/U2  ( .x(\U310_3_/n2 ), .a(\third_ol[3] ) );
    inv_1 \U310_3_/U3  ( .x(\U310_3_/n3 ), .a(\second_ol[3] ) );
    inv_1 \U310_3_/U4  ( .x(\U310_3_/n4 ), .a(\first_ol[3] ) );
    inv_4 \U310_3_/U5  ( .x(ol[3]), .a(\U310_3_/n5 ) );
    and4_2 \U310_4_/U24  ( .x(\U310_4_/n5 ), .a(\U310_4_/n1 ), .b(\U310_4_/n2 
        ), .c(\U310_4_/n3 ), .d(\U310_4_/n4 ) );
    inv_1 \U310_4_/U1  ( .x(\U310_4_/n1 ), .a(\fourth_ol[4] ) );
    inv_1 \U310_4_/U2  ( .x(\U310_4_/n2 ), .a(\third_ol[4] ) );
    inv_1 \U310_4_/U3  ( .x(\U310_4_/n3 ), .a(\second_ol[4] ) );
    inv_1 \U310_4_/U4  ( .x(\U310_4_/n4 ), .a(\first_ol[4] ) );
    inv_4 \U310_4_/U5  ( .x(ol[4]), .a(\U310_4_/n5 ) );
    and4_2 \U310_5_/U24  ( .x(\U310_5_/n5 ), .a(\U310_5_/n1 ), .b(\U310_5_/n2 
        ), .c(\U310_5_/n3 ), .d(\U310_5_/n4 ) );
    inv_1 \U310_5_/U1  ( .x(\U310_5_/n1 ), .a(\fourth_ol[5] ) );
    inv_1 \U310_5_/U2  ( .x(\U310_5_/n2 ), .a(\third_ol[5] ) );
    inv_1 \U310_5_/U3  ( .x(\U310_5_/n3 ), .a(\second_ol[5] ) );
    inv_1 \U310_5_/U4  ( .x(\U310_5_/n4 ), .a(\first_ol[5] ) );
    inv_4 \U310_5_/U5  ( .x(ol[5]), .a(\U310_5_/n5 ) );
    and4_2 \U310_6_/U24  ( .x(\U310_6_/n5 ), .a(\U310_6_/n1 ), .b(\U310_6_/n2 
        ), .c(\U310_6_/n3 ), .d(\U310_6_/n4 ) );
    inv_1 \U310_6_/U1  ( .x(\U310_6_/n1 ), .a(\fourth_ol[6] ) );
    inv_1 \U310_6_/U2  ( .x(\U310_6_/n2 ), .a(\third_ol[6] ) );
    inv_1 \U310_6_/U3  ( .x(\U310_6_/n3 ), .a(\second_ol[6] ) );
    inv_1 \U310_6_/U4  ( .x(\U310_6_/n4 ), .a(\first_ol[6] ) );
    inv_4 \U310_6_/U5  ( .x(ol[6]), .a(\U310_6_/n5 ) );
    and4_2 \U310_7_/U24  ( .x(\U310_7_/n5 ), .a(\U310_7_/n1 ), .b(\U310_7_/n2 
        ), .c(\U310_7_/n3 ), .d(\U310_7_/n4 ) );
    inv_1 \U310_7_/U1  ( .x(\U310_7_/n1 ), .a(\fourth_ol[7] ) );
    inv_1 \U310_7_/U2  ( .x(\U310_7_/n2 ), .a(\third_ol[7] ) );
    inv_1 \U310_7_/U3  ( .x(\U310_7_/n3 ), .a(\second_ol[7] ) );
    inv_1 \U310_7_/U4  ( .x(\U310_7_/n4 ), .a(\first_ol[7] ) );
    inv_4 \U310_7_/U5  ( .x(ol[7]), .a(\U310_7_/n5 ) );
endmodule


module chain_selement_ga_64 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_trhdr_1 ( chainff_ack, chainh, chainl, eop, hdrack, normal_ack, 
    notify_ack, read_req, routereq, chain_ff_h, chainack, chainff_l, eopack, 
    err, nReset, normal_response, notify_accept, notify_defer, rcol_h, rcol_l, 
    read_ack, rnw_h, rnw_l, routeack, rsize_h, rsize_l, rtag_h, rtag_l );
output [7:0] chainh;
output [7:0] chainl;
input  [7:0] chain_ff_h;
input  [7:0] chainff_l;
input  [1:0] err;
input  [2:0] rcol_h;
input  [2:0] rcol_l;
input  [1:0] rsize_h;
input  [1:0] rsize_l;
input  [4:0] rtag_h;
input  [4:0] rtag_l;
input  chainack, eopack, nReset, normal_response, notify_accept, notify_defer, 
    read_ack, rnw_h, rnw_l, routeack;
output chainff_ack, eop, hdrack, normal_ack, notify_ack, read_req, routereq;
    wire \net334[0] , \net334[1] , \net334[2] , \net334[4] , \net334[6] , 
        \net334[7] , \net413[0] , \net413[1] , \net413[2] , \net413[3] , 
        \net413[4] , \net413[5] , \net413[6] , \net413[7] , \net413[8] , 
        \net413[9] , \net413[10] , \net413[11] , \net413[12] , \net413[13] , 
        \net413[14] , \net413[15] , \net284[0] , \net284[1] , \net284[2] , 
        \net284[3] , \net284[4] , \net284[5] , \net284[6] , \net284[7] , 
        \net288[0] , \net288[1] , \net288[2] , \net288[3] , \net288[4] , 
        \net288[5] , \net288[6] , \net288[7] , \net343[0] , \net343[1] , 
        \net343[2] , \net343[3] , \net343[5] , \net343[6] , \net343[7] , 
        \hdr[17] , \hdr[16] , \hdr[1] , \hdr[0] , \drive_h[1] , \drive_h[0] , 
        \drive_l[1] , \drive_l[0] , done_write, dowrite, done_eop, ctrl_cd, 
        done_read, done_hdr, done_defer, net321, net362, net359, done_accept, 
        net332, net337, net340, done_pl, net364, donotify, net383, net0230, 
        net407, \U319/U21/U1/loop , \U323/U21/U1/loop , \U320/U21/U1/loop , 
        \U321/U21/U1/loop , \U322/U21/U1/loop , \U311/U28/Z , \U311/U32/Z , 
        \U311/U20/Z , \U311/U29/Z , \U311/U25/Z , \U311/U33/Z , \U311/U21/Z , 
        \U311/U26/Z , \U311/U34/Z , \U311/U30/Z , \U311/U19/Z , \U311/U27/Z , 
        \U311/U35/Z , \U311/U31/Z , \U311/nz[0] , \U311/nz[1] , \U311/x[1] , 
        \U311/y[3] , \U311/y[2] , \U311/x[7] , \U311/x[6] , \U311/x[4] , 
        \U311/y[1] , \U311/x[3] , \U311/x[2] , \U311/y[0] , \U311/x[5] , 
        \U311/x[0] , \U151/Z , \U210/naa , \U210/bdone , \U210/net3 , 
        \U210/drivemonitor , \U210/net2 , \U210/U1702/Z , \I0/naa , \I0/bdone , 
        \I0/net3 , \I0/drivemonitor , \I0/net2 , \I0/U1702/Z ;
    chain_selement_ga_64 U215 ( .Aa(done_eop), .Br(eop), .Ar(done_pl), .Ba(
        eopack) );
    nor2_1 \U308_0_/U5  ( .x(\net413[15] ), .a(\hdr[16] ), .b(\hdr[0] ) );
    nor2_1 \U308_1_/U5  ( .x(\net413[14] ), .a(\hdr[17] ), .b(\hdr[1] ) );
    nor2_1 \U308_2_/U5  ( .x(\net413[13] ), .a(1'b0), .b(routereq) );
    nor2_1 \U308_3_/U5  ( .x(\net413[12] ), .a(routereq), .b(1'b0) );
    nor2_1 \U308_4_/U5  ( .x(\net413[11] ), .a(1'b0), .b(routereq) );
    nor2_1 \U308_5_/U5  ( .x(\net413[10] ), .a(rnw_h), .b(rnw_l) );
    nor2_1 \U308_6_/U5  ( .x(\net413[9] ), .a(rsize_h[0]), .b(rsize_l[0]) );
    nor2_1 \U308_7_/U5  ( .x(\net413[8] ), .a(rsize_h[1]), .b(rsize_l[1]) );
    nor2_1 \U308_8_/U5  ( .x(\net413[7] ), .a(rtag_h[0]), .b(rtag_l[0]) );
    nor2_1 \U308_9_/U5  ( .x(\net413[6] ), .a(rtag_h[1]), .b(rtag_l[1]) );
    nor2_1 \U308_10_/U5  ( .x(\net413[5] ), .a(rtag_h[2]), .b(rtag_l[2]) );
    nor2_1 \U308_11_/U5  ( .x(\net413[4] ), .a(rtag_h[3]), .b(rtag_l[3]) );
    nor2_1 \U308_12_/U5  ( .x(\net413[3] ), .a(rtag_h[4]), .b(rtag_l[4]) );
    nor2_1 \U308_13_/U5  ( .x(\net413[2] ), .a(rcol_h[0]), .b(rcol_l[0]) );
    nor2_1 \U308_14_/U5  ( .x(\net413[1] ), .a(rcol_h[1]), .b(rcol_l[1]) );
    nor2_1 \U308_15_/U5  ( .x(\net413[0] ), .a(rcol_h[2]), .b(rcol_l[2]) );
    or3_1 \U257/U12  ( .x(net364), .a(donotify), .b(dowrite), .c(read_ack) );
    or3_1 \U297/U12  ( .x(net383), .a(done_defer), .b(done_write), .c(
        done_read) );
    and2_2 \U237/U8  ( .x(\hdr[1] ), .a(nReset), .b(normal_response) );
    and2_1 \U307_0_/U8  ( .x(\net343[7] ), .a(\drive_l[0] ), .b(\hdr[0] ) );
    and2_1 \U307_1_/U8  ( .x(\net343[6] ), .a(\drive_l[0] ), .b(\hdr[1] ) );
    and2_1 \U307_2_/U8  ( .x(\net343[5] ), .a(\drive_l[0] ), .b(routereq) );
    and2_1 \U307_4_/U8  ( .x(\net343[3] ), .a(\drive_l[0] ), .b(routereq) );
    and2_1 \U307_5_/U8  ( .x(\net343[2] ), .a(\drive_l[0] ), .b(rnw_l) );
    and2_1 \U307_6_/U8  ( .x(\net343[1] ), .a(\drive_l[0] ), .b(rsize_l[0]) );
    and2_1 \U307_7_/U8  ( .x(\net343[0] ), .a(\drive_l[0] ), .b(rsize_l[1]) );
    and2_1 \U235/U8  ( .x(net340), .a(err[1]), .b(nReset) );
    and2_1 \U236/U8  ( .x(net337), .a(nReset), .b(err[0]) );
    and2_1 \U306_0_/U8  ( .x(\net334[7] ), .a(\hdr[16] ), .b(\drive_l[1] ) );
    and2_1 \U306_1_/U8  ( .x(\net334[6] ), .a(\hdr[17] ), .b(\drive_l[1] ) );
    and2_1 \U306_3_/U8  ( .x(\net334[4] ), .a(routereq), .b(\drive_l[1] ) );
    and2_1 \U306_5_/U8  ( .x(\net334[2] ), .a(rnw_h), .b(\drive_l[1] ) );
    and2_1 \U306_6_/U8  ( .x(\net334[1] ), .a(rsize_h[0]), .b(\drive_l[1] ) );
    and2_1 \U306_7_/U8  ( .x(\net334[0] ), .a(rsize_h[1]), .b(\drive_l[1] ) );
    and2_1 \I1_0_/U8  ( .x(\net284[7] ), .a(rtag_h[0]), .b(\drive_h[1] ) );
    and2_1 \I1_1_/U8  ( .x(\net284[6] ), .a(rtag_h[1]), .b(\drive_h[1] ) );
    and2_1 \I1_2_/U8  ( .x(\net284[5] ), .a(rtag_h[2]), .b(\drive_h[1] ) );
    and2_1 \I1_3_/U8  ( .x(\net284[4] ), .a(rtag_h[3]), .b(\drive_h[1] ) );
    and2_1 \I1_4_/U8  ( .x(\net284[3] ), .a(rtag_h[4]), .b(\drive_h[1] ) );
    and2_1 \I1_5_/U8  ( .x(\net284[2] ), .a(rcol_h[0]), .b(\drive_h[1] ) );
    and2_1 \I1_6_/U8  ( .x(\net284[1] ), .a(rcol_h[1]), .b(\drive_h[1] ) );
    and2_1 \I1_7_/U8  ( .x(\net284[0] ), .a(rcol_h[2]), .b(\drive_h[1] ) );
    and2_1 \I2_0_/U8  ( .x(\net288[7] ), .a(\drive_h[0] ), .b(rtag_l[0]) );
    and2_1 \I2_1_/U8  ( .x(\net288[6] ), .a(\drive_h[0] ), .b(rtag_l[1]) );
    and2_1 \I2_2_/U8  ( .x(\net288[5] ), .a(\drive_h[0] ), .b(rtag_l[2]) );
    and2_1 \I2_3_/U8  ( .x(\net288[4] ), .a(\drive_h[0] ), .b(rtag_l[3]) );
    and2_1 \I2_4_/U8  ( .x(\net288[3] ), .a(\drive_h[0] ), .b(rtag_l[4]) );
    and2_1 \I2_5_/U8  ( .x(\net288[2] ), .a(\drive_h[0] ), .b(rcol_l[0]) );
    and2_1 \I2_6_/U8  ( .x(\net288[1] ), .a(\drive_h[0] ), .b(rcol_l[1]) );
    and2_1 \I2_7_/U8  ( .x(\net288[0] ), .a(\drive_h[0] ), .b(rcol_l[2]) );
    inv_1 \U318/U3  ( .x(net332), .a(routereq) );
    or2_4 \U255/U12  ( .x(notify_ack), .a(done_accept), .b(done_defer) );
    or2_4 \U228/U12  ( .x(\hdr[17] ), .a(notify_defer), .b(notify_accept) );
    or2_4 \U204/U12  ( .x(net321), .a(net359), .b(net362) );
    or2_4 \U221/U12  ( .x(\hdr[16] ), .a(net359), .b(notify_defer) );
    or2_4 \U252/U12  ( .x(normal_ack), .a(done_write), .b(done_read) );
    or2_4 \U280/U12  ( .x(\hdr[0] ), .a(net362), .b(notify_accept) );
    or2_4 \U317/U12  ( .x(routereq), .a(\hdr[17] ), .b(net321) );
    or3_4 \U309_0_/U12  ( .x(chainh[0]), .a(\net334[7] ), .b(\net284[7] ), .c(
        chain_ff_h[0]) );
    or3_4 \U309_1_/U12  ( .x(chainh[1]), .a(\net334[6] ), .b(\net284[6] ), .c(
        chain_ff_h[1]) );
    or3_4 \U309_3_/U12  ( .x(chainh[3]), .a(\net334[4] ), .b(\net284[4] ), .c(
        chain_ff_h[3]) );
    or3_4 \U309_5_/U12  ( .x(chainh[5]), .a(\net334[2] ), .b(\net284[2] ), .c(
        chain_ff_h[5]) );
    or3_4 \U309_6_/U12  ( .x(chainh[6]), .a(\net334[1] ), .b(\net284[1] ), .c(
        chain_ff_h[6]) );
    or3_4 \U309_7_/U12  ( .x(chainh[7]), .a(\net334[0] ), .b(\net284[0] ), .c(
        chain_ff_h[7]) );
    or3_4 \U310_0_/U12  ( .x(chainl[0]), .a(\net343[7] ), .b(\net288[7] ), .c(
        chainff_l[0]) );
    or3_4 \U310_1_/U12  ( .x(chainl[1]), .a(\net343[6] ), .b(\net288[6] ), .c(
        chainff_l[1]) );
    or3_4 \U310_2_/U12  ( .x(chainl[2]), .a(\net343[5] ), .b(\net288[5] ), .c(
        chainff_l[2]) );
    or3_4 \U310_4_/U12  ( .x(chainl[4]), .a(\net343[3] ), .b(\net288[3] ), .c(
        chainff_l[4]) );
    or3_4 \U310_5_/U12  ( .x(chainl[5]), .a(\net343[2] ), .b(\net288[2] ), .c(
        chainff_l[5]) );
    or3_4 \U310_6_/U12  ( .x(chainl[6]), .a(\net343[1] ), .b(\net288[1] ), .c(
        chainff_l[6]) );
    or3_4 \U310_7_/U12  ( .x(chainl[7]), .a(\net343[0] ), .b(\net288[0] ), .c(
        chainff_l[7]) );
    ao222_1 \U311/U37/U18/U1/U1  ( .x(ctrl_cd), .a(\U311/nz[0] ), .b(
        \U311/nz[1] ), .c(\U311/nz[0] ), .d(ctrl_cd), .e(\U311/nz[1] ), .f(
        ctrl_cd) );
    aoi222_1 \U311/U28/U30/U1  ( .x(\U311/x[3] ), .a(\net413[8] ), .b(
        \net413[9] ), .c(\net413[8] ), .d(\U311/U28/Z ), .e(\net413[9] ), .f(
        \U311/U28/Z ) );
    inv_1 \U311/U28/U30/Uinv  ( .x(\U311/U28/Z ), .a(\U311/x[3] ) );
    aoi222_1 \U311/U32/U30/U1  ( .x(\U311/x[0] ), .a(\net413[14] ), .b(
        \net413[15] ), .c(\net413[14] ), .d(\U311/U32/Z ), .e(\net413[15] ), 
        .f(\U311/U32/Z ) );
    inv_1 \U311/U32/U30/Uinv  ( .x(\U311/U32/Z ), .a(\U311/x[0] ) );
    aoi222_1 \U311/U20/U30/U1  ( .x(\U311/x[5] ), .a(\net413[4] ), .b(
        \net413[5] ), .c(\net413[4] ), .d(\U311/U20/Z ), .e(\net413[5] ), .f(
        \U311/U20/Z ) );
    inv_1 \U311/U20/U30/Uinv  ( .x(\U311/U20/Z ), .a(\U311/x[5] ) );
    aoi222_1 \U311/U29/U30/U1  ( .x(\U311/x[2] ), .a(\net413[10] ), .b(
        \net413[11] ), .c(\net413[10] ), .d(\U311/U29/Z ), .e(\net413[11] ), 
        .f(\U311/U29/Z ) );
    inv_1 \U311/U29/U30/Uinv  ( .x(\U311/U29/Z ), .a(\U311/x[2] ) );
    aoi222_1 \U311/U25/U30/U1  ( .x(\U311/x[7] ), .a(\net413[0] ), .b(
        \net413[1] ), .c(\net413[0] ), .d(\U311/U25/Z ), .e(\net413[1] ), .f(
        \U311/U25/Z ) );
    inv_1 \U311/U25/U30/Uinv  ( .x(\U311/U25/Z ), .a(\U311/x[7] ) );
    aoi222_1 \U311/U33/U30/U1  ( .x(\U311/y[0] ), .a(\U311/x[1] ), .b(
        \U311/x[0] ), .c(\U311/x[1] ), .d(\U311/U33/Z ), .e(\U311/x[0] ), .f(
        \U311/U33/Z ) );
    inv_1 \U311/U33/U30/Uinv  ( .x(\U311/U33/Z ), .a(\U311/y[0] ) );
    aoi222_1 \U311/U21/U30/U1  ( .x(\U311/y[2] ), .a(\U311/x[5] ), .b(
        \U311/x[4] ), .c(\U311/x[5] ), .d(\U311/U21/Z ), .e(\U311/x[4] ), .f(
        \U311/U21/Z ) );
    inv_1 \U311/U21/U30/Uinv  ( .x(\U311/U21/Z ), .a(\U311/y[2] ) );
    aoi222_1 \U311/U26/U30/U1  ( .x(\U311/x[6] ), .a(\net413[2] ), .b(
        \net413[3] ), .c(\net413[2] ), .d(\U311/U26/Z ), .e(\net413[3] ), .f(
        \U311/U26/Z ) );
    inv_1 \U311/U26/U30/Uinv  ( .x(\U311/U26/Z ), .a(\U311/x[6] ) );
    aoi222_1 \U311/U34/U30/U1  ( .x(\U311/nz[0] ), .a(\U311/y[1] ), .b(
        \U311/y[0] ), .c(\U311/y[1] ), .d(\U311/U34/Z ), .e(\U311/y[0] ), .f(
        \U311/U34/Z ) );
    inv_1 \U311/U34/U30/Uinv  ( .x(\U311/U34/Z ), .a(\U311/nz[0] ) );
    aoi222_1 \U311/U30/U30/U1  ( .x(\U311/y[1] ), .a(\U311/x[3] ), .b(
        \U311/x[2] ), .c(\U311/x[3] ), .d(\U311/U30/Z ), .e(\U311/x[2] ), .f(
        \U311/U30/Z ) );
    inv_1 \U311/U30/U30/Uinv  ( .x(\U311/U30/Z ), .a(\U311/y[1] ) );
    aoi222_1 \U311/U19/U30/U1  ( .x(\U311/x[4] ), .a(\net413[6] ), .b(
        \net413[7] ), .c(\net413[6] ), .d(\U311/U19/Z ), .e(\net413[7] ), .f(
        \U311/U19/Z ) );
    inv_1 \U311/U19/U30/Uinv  ( .x(\U311/U19/Z ), .a(\U311/x[4] ) );
    aoi222_1 \U311/U27/U30/U1  ( .x(\U311/y[3] ), .a(\U311/x[7] ), .b(
        \U311/x[6] ), .c(\U311/x[7] ), .d(\U311/U27/Z ), .e(\U311/x[6] ), .f(
        \U311/U27/Z ) );
    inv_1 \U311/U27/U30/Uinv  ( .x(\U311/U27/Z ), .a(\U311/y[3] ) );
    aoi222_1 \U311/U35/U30/U1  ( .x(\U311/nz[1] ), .a(\U311/y[3] ), .b(
        \U311/y[2] ), .c(\U311/y[3] ), .d(\U311/U35/Z ), .e(\U311/y[2] ), .f(
        \U311/U35/Z ) );
    inv_1 \U311/U35/U30/Uinv  ( .x(\U311/U35/Z ), .a(\U311/nz[1] ) );
    aoi222_1 \U311/U31/U30/U1  ( .x(\U311/x[1] ), .a(\net413[12] ), .b(
        \net413[13] ), .c(\net413[12] ), .d(\U311/U31/Z ), .e(\net413[13] ), 
        .f(\U311/U31/Z ) );
    inv_1 \U311/U31/U30/Uinv  ( .x(\U311/U31/Z ), .a(\U311/x[1] ) );
    aoi21_1 \U151/U30/U1/U1  ( .x(net407), .a(\U151/Z ), .b(chainff_ack), .c(
        net332) );
    inv_1 \U151/U30/U1/U2  ( .x(\U151/Z ), .a(net407) );
    ao222_1 \U324/U18/U1/U1  ( .x(hdrack), .a(ctrl_cd), .b(net383), .c(ctrl_cd
        ), .d(hdrack), .e(net383), .f(hdrack) );
    ao222_1 \U244/U18/U1/U1  ( .x(donotify), .a(done_hdr), .b(\hdr[17] ), .c(
        done_hdr), .d(donotify), .e(\hdr[17] ), .f(donotify) );
    ao222_1 \U260/U18/U1/U1  ( .x(net362), .a(net337), .b(\hdr[1] ), .c(net337
        ), .d(net362), .e(\hdr[1] ), .f(net362) );
    ao222_1 \U296/U18/U1/U1  ( .x(done_accept), .a(done_eop), .b(notify_accept
        ), .c(done_eop), .d(done_accept), .e(notify_accept), .f(done_accept)
         );
    ao222_1 \U261/U18/U1/U1  ( .x(net359), .a(net340), .b(\hdr[1] ), .c(net340
        ), .d(net359), .e(\hdr[1] ), .f(net359) );
    ao222_1 \U316/U18/U1/U1  ( .x(done_pl), .a(net364), .b(routeack), .c(
        net364), .d(done_pl), .e(routeack), .f(done_pl) );
    ao31_1 \U319/U21/U1/aoi  ( .x(\U319/U21/U1/loop ), .a(\hdr[1] ), .b(
        done_hdr), .c(rnw_h), .d(read_req) );
    oa21_1 \U319/U21/U1/outGate  ( .x(read_req), .a(\hdr[1] ), .b(done_hdr), 
        .c(\U319/U21/U1/loop ) );
    ao31_1 \U323/U21/U1/aoi  ( .x(\U323/U21/U1/loop ), .a(done_eop), .b(
        notify_defer), .c(ctrl_cd), .d(done_defer) );
    oa21_1 \U323/U21/U1/outGate  ( .x(done_defer), .a(done_eop), .b(
        notify_defer), .c(\U323/U21/U1/loop ) );
    ao31_1 \U320/U21/U1/aoi  ( .x(\U320/U21/U1/loop ), .a(\hdr[1] ), .b(
        done_hdr), .c(rnw_l), .d(dowrite) );
    oa21_1 \U320/U21/U1/outGate  ( .x(dowrite), .a(\hdr[1] ), .b(done_hdr), 
        .c(\U320/U21/U1/loop ) );
    ao31_1 \U321/U21/U1/aoi  ( .x(\U321/U21/U1/loop ), .a(read_req), .b(
        done_eop), .c(ctrl_cd), .d(done_read) );
    oa21_1 \U321/U21/U1/outGate  ( .x(done_read), .a(read_req), .b(done_eop), 
        .c(\U321/U21/U1/loop ) );
    ao31_1 \U322/U21/U1/aoi  ( .x(\U322/U21/U1/loop ), .a(dowrite), .b(
        done_eop), .c(ctrl_cd), .d(done_write) );
    oa21_1 \U322/U21/U1/outGate  ( .x(done_write), .a(dowrite), .b(done_eop), 
        .c(\U322/U21/U1/loop ) );
    nor2_2 \U210/U1703/U6  ( .x(done_hdr), .a(\U210/drivemonitor ), .b(
        \U210/naa ) );
    inv_2 \U210/U1699/U3  ( .x(\U210/net2 ), .a(\U210/net3 ) );
    and2_4 \U210/U2_0_/U8  ( .x(\drive_l[0] ), .a(net0230), .b(\U210/net2 ) );
    and2_4 \U210/U2_1_/U8  ( .x(\drive_l[1] ), .a(net0230), .b(\U210/net2 ) );
    inv_1 \U210/U1701/U3  ( .x(\U210/naa ), .a(\U210/bdone ) );
    ao222_1 \U210/U13/U18/U1/U1  ( .x(\U210/drivemonitor ), .a(\drive_l[1] ), 
        .b(\drive_l[0] ), .c(\drive_l[1] ), .d(\U210/drivemonitor ), .e(
        \drive_l[0] ), .f(\U210/drivemonitor ) );
    aoi21_1 \U210/U1702/U30/U1/U1  ( .x(\U210/bdone ), .a(\U210/U1702/Z ), .b(
        chainff_ack), .c(\U210/net2 ) );
    inv_1 \U210/U1702/U30/U1/U2  ( .x(\U210/U1702/Z ), .a(\U210/bdone ) );
    ao23_1 \U210/U1693/U21/U1/U1  ( .x(\U210/net3 ), .a(net0230), .b(
        \U210/net3 ), .c(net0230), .d(\U210/drivemonitor ), .e(chainff_ack) );
    nor2_2 \I0/U1703/U6  ( .x(net0230), .a(\I0/drivemonitor ), .b(\I0/naa ) );
    inv_2 \I0/U1699/U3  ( .x(\I0/net2 ), .a(\I0/net3 ) );
    and2_4 \I0/U2_0_/U8  ( .x(\drive_h[0] ), .a(net407), .b(\I0/net2 ) );
    and2_4 \I0/U2_1_/U8  ( .x(\drive_h[1] ), .a(net407), .b(\I0/net2 ) );
    inv_1 \I0/U1701/U3  ( .x(\I0/naa ), .a(\I0/bdone ) );
    ao222_1 \I0/U13/U18/U1/U1  ( .x(\I0/drivemonitor ), .a(\drive_h[1] ), .b(
        \drive_h[0] ), .c(\drive_h[1] ), .d(\I0/drivemonitor ), .e(
        \drive_h[0] ), .f(\I0/drivemonitor ) );
    aoi21_1 \I0/U1702/U30/U1/U1  ( .x(\I0/bdone ), .a(\I0/U1702/Z ), .b(
        chainff_ack), .c(\I0/net2 ) );
    inv_1 \I0/U1702/U30/U1/U2  ( .x(\I0/U1702/Z ), .a(\I0/bdone ) );
    ao23_1 \I0/U1693/U21/U1/U1  ( .x(\I0/net3 ), .a(net407), .b(\I0/net3 ), 
        .c(net407), .d(\I0/drivemonitor ), .e(chainff_ack) );
    buf_3 U1 ( .x(chainff_ack), .a(chainack) );
    or2_1 U2 ( .x(chainh[4]), .a(chain_ff_h[4]), .b(\net284[3] ) );
    or2_1 U3 ( .x(chainh[2]), .a(chain_ff_h[2]), .b(\net284[5] ) );
    or2_1 U4 ( .x(chainl[3]), .a(chainff_l[3]), .b(\net288[4] ) );
endmodule


module chain_tchdr_1 ( addr_req, col_h, col_l, itag_h, itag_l, lock, ncback, 
    neop, pred, pullcd, reset, rnw_h, rnw_l, seq, size_h, size_l, write_req, 
    chwh, chwl, addr_ack, addr_pull, nReset, nack, write_ack, write_pull );
output [2:0] col_h;
output [2:0] col_l;
output [4:0] itag_h;
output [4:0] itag_l;
output [1:0] lock;
output [1:0] pred;
output [1:0] seq;
output [1:0] size_h;
output [1:0] size_l;
input  [7:0] chwh;
input  [7:0] chwl;
input  addr_ack, addr_pull, nReset, nack, write_ack, write_pull;
output addr_req, ncback, neop, pullcd, reset, rnw_h, rnw_l, write_req;
    wire \ncd[7] , \ncd[6] , \ncd[5] , \ncd[4] , \ncd[3] , \ncd[2] , \ncd[1] , 
        \ncd[0] , net88, receive, pullcdwk, read, net83, ack, net94, n9, 
        \U1664/U28/Z , \U1664/U32/Z , \U1664/U29/Z , \U1664/U33/Z , 
        \U1664/U30/Z , \U1664/U31/Z , \U1664/U37/Z , \U473/Z , \U1664/y[0] , 
        \U1664/y[1] , \U1664/x[1] , \U1664/x[3] , \U1664/x[2] , \U1664/x[0] , 
        \hdr_hld/oh[4] , \hdr_hld/oh[3] , \hdr_hld/ol[4] , \hdr_hld/ol[3] , 
        \hdr_hld/net20 , \hdr_hld/net33 , \hdr_hld/net32 , 
        \hdr_hld/low/drivel , \hdr_hld/low/driveh , \hdr_hld/low/localcd , 
        \hdr_hld/low/ncd[7] , \hdr_hld/low/ncd[6] , \hdr_hld/low/ncd[5] , 
        \hdr_hld/low/ncd[4] , \hdr_hld/low/ncd[3] , \hdr_hld/low/ncd[2] , 
        \hdr_hld/low/ncd[1] , \hdr_hld/low/ncd[0] , \hdr_hld/low/ba , 
        \hdr_hld/low/latch , \hdr_hld/low/acb , \hdr_hld/low/ctrlack_internal , 
        \hdr_hld/low/nlocalcd , \hdr_hld/low/U4/U28/U1/clr , 
        \hdr_hld/low/U4/U28/U1/set , \hdr_hld/low/U1/Z , 
        \hdr_hld/low/U1664/y[0] , \hdr_hld/low/U1664/y[1] , 
        \hdr_hld/low/U1664/x[1] , \hdr_hld/low/U1664/x[3] , 
        \hdr_hld/low/U1664/x[2] , \hdr_hld/low/U1664/x[0] , 
        \hdr_hld/low/U1664/U28/Z , \hdr_hld/low/U1664/U32/Z , 
        \hdr_hld/low/U1664/U29/Z , \hdr_hld/low/U1664/U33/Z , 
        \hdr_hld/low/U1664/U30/Z , \hdr_hld/low/U1664/U31/Z , 
        \hdr_hld/low/U1664/U37/Z , \hdr_hld/low/U1669/nr , 
        \hdr_hld/low/U1669/nd , \hdr_hld/low/U1669/n2 , \hdr_hld/high/drivel , 
        \hdr_hld/high/driveh , \hdr_hld/high/localcd , \hdr_hld/high/ncd[7] , 
        \hdr_hld/high/ncd[6] , \hdr_hld/high/ncd[5] , \hdr_hld/high/ncd[4] , 
        \hdr_hld/high/ncd[3] , \hdr_hld/high/ncd[2] , \hdr_hld/high/ncd[1] , 
        \hdr_hld/high/ncd[0] , \hdr_hld/high/ba , \hdr_hld/high/latch , 
        \hdr_hld/high/acb , \hdr_hld/high/ctrlack_internal , 
        \hdr_hld/high/nlocalcd , \hdr_hld/high/U4/U28/U1/clr , 
        \hdr_hld/high/U4/U28/U1/set , \hdr_hld/high/U1/Z , 
        \hdr_hld/high/U1664/y[0] , \hdr_hld/high/U1664/y[1] , 
        \hdr_hld/high/U1664/x[1] , \hdr_hld/high/U1664/x[3] , 
        \hdr_hld/high/U1664/x[2] , \hdr_hld/high/U1664/x[0] , 
        \hdr_hld/high/U1664/U28/Z , \hdr_hld/high/U1664/U32/Z , 
        \hdr_hld/high/U1664/U29/Z , \hdr_hld/high/U1664/U33/Z , 
        \hdr_hld/high/U1664/U30/Z , \hdr_hld/high/U1664/U31/Z , 
        \hdr_hld/high/U1664/U37/Z , \hdr_hld/high/U1669/nr , 
        \hdr_hld/high/U1669/nd , \hdr_hld/high/U1669/n2 , n1, n2, n3, n4, n5, 
        n6, n7;
    buf_1 U262 ( .x(n9), .a(pullcdwk) );
    or3_2 \U1668/U12  ( .x(ncback), .a(net94), .b(addr_pull), .c(write_pull)
         );
    inv_1 \I0/U3  ( .x(net94), .a(net88) );
    nor2_1 \U514_0_/U5  ( .x(\ncd[0] ), .a(chwh[0]), .b(chwl[0]) );
    nor2_1 \U514_1_/U5  ( .x(\ncd[1] ), .a(chwh[1]), .b(chwl[1]) );
    nor2_1 \U514_2_/U5  ( .x(\ncd[2] ), .a(chwh[2]), .b(chwl[2]) );
    nor2_1 \U514_3_/U5  ( .x(\ncd[3] ), .a(chwh[3]), .b(chwl[3]) );
    nor2_1 \U514_4_/U5  ( .x(\ncd[4] ), .a(chwh[4]), .b(chwl[4]) );
    nor2_1 \U514_5_/U5  ( .x(\ncd[5] ), .a(chwh[5]), .b(chwl[5]) );
    nor2_1 \U514_6_/U5  ( .x(\ncd[6] ), .a(chwh[6]), .b(chwl[6]) );
    nor2_1 \U514_7_/U5  ( .x(\ncd[7] ), .a(chwh[7]), .b(chwl[7]) );
    nor2_1 \U1669/U5  ( .x(neop), .a(read), .b(write_ack) );
    nand2_1 \U303/U5  ( .x(ack), .a(nack), .b(nReset) );
    nand2_1 \U1670/U5  ( .x(net83), .a(neop), .b(nReset) );
    ao222_1 \U47/U18/U1/U1  ( .x(read), .a(addr_ack), .b(rnw_h), .c(addr_ack), 
        .d(read), .e(rnw_h), .f(read) );
    ao222_1 \U48/U18/U1/U1  ( .x(write_req), .a(rnw_l), .b(addr_ack), .c(rnw_l
        ), .d(write_req), .e(addr_ack), .f(write_req) );
    aoi222_1 \U1664/U28/U30/U1  ( .x(\U1664/x[3] ), .a(\ncd[7] ), .b(\ncd[6] ), 
        .c(\ncd[7] ), .d(\U1664/U28/Z ), .e(\ncd[6] ), .f(\U1664/U28/Z ) );
    inv_1 \U1664/U28/U30/Uinv  ( .x(\U1664/U28/Z ), .a(\U1664/x[3] ) );
    aoi222_1 \U1664/U32/U30/U1  ( .x(\U1664/x[0] ), .a(\ncd[1] ), .b(\ncd[0] ), 
        .c(\ncd[1] ), .d(\U1664/U32/Z ), .e(\ncd[0] ), .f(\U1664/U32/Z ) );
    inv_1 \U1664/U32/U30/Uinv  ( .x(\U1664/U32/Z ), .a(\U1664/x[0] ) );
    aoi222_1 \U1664/U29/U30/U1  ( .x(\U1664/x[2] ), .a(\ncd[5] ), .b(\ncd[4] ), 
        .c(\ncd[5] ), .d(\U1664/U29/Z ), .e(\ncd[4] ), .f(\U1664/U29/Z ) );
    inv_1 \U1664/U29/U30/Uinv  ( .x(\U1664/U29/Z ), .a(\U1664/x[2] ) );
    aoi222_1 \U1664/U33/U30/U1  ( .x(\U1664/y[0] ), .a(\U1664/x[1] ), .b(
        \U1664/x[0] ), .c(\U1664/x[1] ), .d(\U1664/U33/Z ), .e(\U1664/x[0] ), 
        .f(\U1664/U33/Z ) );
    inv_1 \U1664/U33/U30/Uinv  ( .x(\U1664/U33/Z ), .a(\U1664/y[0] ) );
    aoi222_1 \U1664/U30/U30/U1  ( .x(\U1664/y[1] ), .a(\U1664/x[3] ), .b(
        \U1664/x[2] ), .c(\U1664/x[3] ), .d(\U1664/U30/Z ), .e(\U1664/x[2] ), 
        .f(\U1664/U30/Z ) );
    inv_1 \U1664/U30/U30/Uinv  ( .x(\U1664/U30/Z ), .a(\U1664/y[1] ) );
    aoi222_1 \U1664/U31/U30/U1  ( .x(\U1664/x[1] ), .a(\ncd[3] ), .b(\ncd[2] ), 
        .c(\ncd[3] ), .d(\U1664/U31/Z ), .e(\ncd[2] ), .f(\U1664/U31/Z ) );
    inv_1 \U1664/U31/U30/Uinv  ( .x(\U1664/U31/Z ), .a(\U1664/x[1] ) );
    aoi222_1 \U1664/U37/U30/U1  ( .x(pullcdwk), .a(\U1664/y[0] ), .b(
        \U1664/y[1] ), .c(\U1664/y[0] ), .d(\U1664/U37/Z ), .e(\U1664/y[1] ), 
        .f(\U1664/U37/Z ) );
    inv_1 \U1664/U37/U30/Uinv  ( .x(\U1664/U37/Z ), .a(pullcdwk) );
    aoi222_1 \U473/U30/U1  ( .x(receive), .a(net83), .b(ack), .c(net83), .d(
        \U473/Z ), .e(ack), .f(\U473/Z ) );
    inv_1 \U473/U30/Uinv  ( .x(\U473/Z ), .a(receive) );
    nor2_1 \hdr_hld/U3/U5  ( .x(net88), .a(\hdr_hld/net32 ), .b(
        \hdr_hld/net33 ) );
    buf_2 \hdr_hld/low/U1653  ( .x(\hdr_hld/low/latch ), .a(\hdr_hld/net32 )
         );
    nor2_1 \hdr_hld/low/U264/U5  ( .x(\hdr_hld/low/nlocalcd ), .a(reset), .b(
        \hdr_hld/low/localcd ) );
    nor2_1 \hdr_hld/low/U1659_0_/U5  ( .x(\hdr_hld/low/ncd[0] ), .a(seq[0]), 
        .b(seq[1]) );
    nor2_1 \hdr_hld/low/U1659_1_/U5  ( .x(\hdr_hld/low/ncd[1] ), .a(pred[0]), 
        .b(pred[1]) );
    nor2_1 \hdr_hld/low/U1659_2_/U5  ( .x(\hdr_hld/low/ncd[2] ), .a(lock[0]), 
        .b(lock[1]) );
    nor2_1 \hdr_hld/low/U1659_3_/U5  ( .x(\hdr_hld/low/ncd[3] ), .a(
        \hdr_hld/ol[3] ), .b(\hdr_hld/oh[3] ) );
    nor2_1 \hdr_hld/low/U1659_4_/U5  ( .x(\hdr_hld/low/ncd[4] ), .a(
        \hdr_hld/ol[4] ), .b(\hdr_hld/oh[4] ) );
    nor2_1 \hdr_hld/low/U1659_5_/U5  ( .x(\hdr_hld/low/ncd[5] ), .a(rnw_l), 
        .b(rnw_h) );
    nor2_1 \hdr_hld/low/U1659_6_/U5  ( .x(\hdr_hld/low/ncd[6] ), .a(size_l[0]), 
        .b(size_h[0]) );
    nor2_1 \hdr_hld/low/U1659_7_/U5  ( .x(\hdr_hld/low/ncd[7] ), .a(size_l[1]), 
        .b(size_h[1]) );
    nor2_1 \hdr_hld/low/U3/U5  ( .x(\hdr_hld/low/ctrlack_internal ), .a(
        \hdr_hld/low/acb ), .b(\hdr_hld/low/ba ) );
    buf_2 \hdr_hld/low/U1665/U7  ( .x(\hdr_hld/low/driveh ), .a(
        \hdr_hld/net20 ) );
    buf_2 \hdr_hld/low/U1666/U7  ( .x(\hdr_hld/low/drivel ), .a(
        \hdr_hld/net20 ) );
    ao23_1 \hdr_hld/low/U1658_0_/U21/U1/U1  ( .x(seq[0]), .a(n2), .b(seq[0]), 
        .c(\hdr_hld/low/drivel ), .d(chwl[0]), .e(n3) );
    ao23_1 \hdr_hld/low/U1658_1_/U21/U1/U1  ( .x(pred[0]), .a(n1), .b(pred[0]), 
        .c(\hdr_hld/low/drivel ), .d(chwl[1]), .e(n3) );
    ao23_1 \hdr_hld/low/U1658_2_/U21/U1/U1  ( .x(lock[0]), .a(n1), .b(lock[0]), 
        .c(\hdr_hld/low/driveh ), .d(chwl[2]), .e(n3) );
    ao23_1 \hdr_hld/low/U1658_3_/U21/U1/U1  ( .x(\hdr_hld/ol[3] ), .a(n1), .b(
        \hdr_hld/ol[3] ), .c(\hdr_hld/low/driveh ), .d(chwl[3]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_4_/U21/U1/U1  ( .x(\hdr_hld/ol[4] ), .a(n2), .b(
        \hdr_hld/ol[4] ), .c(\hdr_hld/low/drivel ), .d(chwl[4]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_5_/U21/U1/U1  ( .x(rnw_l), .a(
        \hdr_hld/low/driveh ), .b(rnw_l), .c(\hdr_hld/low/driveh ), .d(chwl[5]
        ), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_6_/U21/U1/U1  ( .x(size_l[0]), .a(
        \hdr_hld/low/drivel ), .b(size_l[0]), .c(n2), .d(chwl[6]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_7_/U21/U1/U1  ( .x(size_l[1]), .a(
        \hdr_hld/low/drivel ), .b(size_l[1]), .c(\hdr_hld/low/drivel ), .d(
        chwl[7]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_0_/U21/U1/U1  ( .x(seq[1]), .a(
        \hdr_hld/low/drivel ), .b(seq[1]), .c(\hdr_hld/low/driveh ), .d(chwh
        [0]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_1_/U21/U1/U1  ( .x(pred[1]), .a(
        \hdr_hld/low/driveh ), .b(pred[1]), .c(n1), .d(chwh[1]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_2_/U21/U1/U1  ( .x(lock[1]), .a(
        \hdr_hld/low/driveh ), .b(lock[1]), .c(n1), .d(chwh[2]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_3_/U21/U1/U1  ( .x(\hdr_hld/oh[3] ), .a(
        \hdr_hld/low/drivel ), .b(\hdr_hld/oh[3] ), .c(n2), .d(chwh[3]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_4_/U21/U1/U1  ( .x(\hdr_hld/oh[4] ), .a(n2), .b(
        \hdr_hld/oh[4] ), .c(n1), .d(chwh[4]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_5_/U21/U1/U1  ( .x(rnw_h), .a(n2), .b(rnw_h), 
        .c(n1), .d(chwh[5]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_6_/U21/U1/U1  ( .x(size_h[0]), .a(n1), .b(size_h
        [0]), .c(n2), .d(chwh[6]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_7_/U21/U1/U1  ( .x(size_h[1]), .a(
        \hdr_hld/low/driveh ), .b(size_h[1]), .c(n2), .d(chwh[7]), .e(
        \hdr_hld/low/latch ) );
    aoai211_1 \hdr_hld/low/U4/U28/U1/U1  ( .x(\hdr_hld/low/U4/U28/U1/clr ), 
        .a(\hdr_hld/net20 ), .b(\hdr_hld/low/acb ), .c(\hdr_hld/low/nlocalcd ), 
        .d(\hdr_hld/net32 ) );
    nand3_1 \hdr_hld/low/U4/U28/U1/U2  ( .x(\hdr_hld/low/U4/U28/U1/set ), .a(
        \hdr_hld/low/nlocalcd ), .b(\hdr_hld/net20 ), .c(\hdr_hld/low/acb ) );
    nand2_2 \hdr_hld/low/U4/U28/U1/U3  ( .x(\hdr_hld/net32 ), .a(
        \hdr_hld/low/U4/U28/U1/clr ), .b(\hdr_hld/low/U4/U28/U1/set ) );
    oai21_1 \hdr_hld/low/U1/U30/U1/U1  ( .x(\hdr_hld/low/acb ), .a(
        \hdr_hld/low/U1/Z ), .b(\hdr_hld/low/ba ), .c(\hdr_hld/net20 ) );
    inv_1 \hdr_hld/low/U1/U30/U1/U2  ( .x(\hdr_hld/low/U1/Z ), .a(
        \hdr_hld/low/acb ) );
    ao222_1 \hdr_hld/low/U5/U18/U1/U1  ( .x(\hdr_hld/low/ba ), .a(
        \hdr_hld/low/latch ), .b(n9), .c(\hdr_hld/low/latch ), .d(
        \hdr_hld/low/ba ), .e(n9), .f(\hdr_hld/low/ba ) );
    aoi222_1 \hdr_hld/low/U1664/U28/U30/U1  ( .x(\hdr_hld/low/U1664/x[3] ), 
        .a(\hdr_hld/low/ncd[7] ), .b(\hdr_hld/low/ncd[6] ), .c(
        \hdr_hld/low/ncd[7] ), .d(\hdr_hld/low/U1664/U28/Z ), .e(
        \hdr_hld/low/ncd[6] ), .f(\hdr_hld/low/U1664/U28/Z ) );
    inv_1 \hdr_hld/low/U1664/U28/U30/Uinv  ( .x(\hdr_hld/low/U1664/U28/Z ), 
        .a(\hdr_hld/low/U1664/x[3] ) );
    aoi222_1 \hdr_hld/low/U1664/U32/U30/U1  ( .x(\hdr_hld/low/U1664/x[0] ), 
        .a(\hdr_hld/low/ncd[1] ), .b(\hdr_hld/low/ncd[0] ), .c(
        \hdr_hld/low/ncd[1] ), .d(\hdr_hld/low/U1664/U32/Z ), .e(
        \hdr_hld/low/ncd[0] ), .f(\hdr_hld/low/U1664/U32/Z ) );
    inv_1 \hdr_hld/low/U1664/U32/U30/Uinv  ( .x(\hdr_hld/low/U1664/U32/Z ), 
        .a(\hdr_hld/low/U1664/x[0] ) );
    aoi222_1 \hdr_hld/low/U1664/U29/U30/U1  ( .x(\hdr_hld/low/U1664/x[2] ), 
        .a(\hdr_hld/low/ncd[5] ), .b(\hdr_hld/low/ncd[4] ), .c(
        \hdr_hld/low/ncd[5] ), .d(\hdr_hld/low/U1664/U29/Z ), .e(
        \hdr_hld/low/ncd[4] ), .f(\hdr_hld/low/U1664/U29/Z ) );
    inv_1 \hdr_hld/low/U1664/U29/U30/Uinv  ( .x(\hdr_hld/low/U1664/U29/Z ), 
        .a(\hdr_hld/low/U1664/x[2] ) );
    aoi222_1 \hdr_hld/low/U1664/U33/U30/U1  ( .x(\hdr_hld/low/U1664/y[0] ), 
        .a(\hdr_hld/low/U1664/x[1] ), .b(\hdr_hld/low/U1664/x[0] ), .c(
        \hdr_hld/low/U1664/x[1] ), .d(\hdr_hld/low/U1664/U33/Z ), .e(
        \hdr_hld/low/U1664/x[0] ), .f(\hdr_hld/low/U1664/U33/Z ) );
    inv_1 \hdr_hld/low/U1664/U33/U30/Uinv  ( .x(\hdr_hld/low/U1664/U33/Z ), 
        .a(\hdr_hld/low/U1664/y[0] ) );
    aoi222_1 \hdr_hld/low/U1664/U30/U30/U1  ( .x(\hdr_hld/low/U1664/y[1] ), 
        .a(\hdr_hld/low/U1664/x[3] ), .b(\hdr_hld/low/U1664/x[2] ), .c(
        \hdr_hld/low/U1664/x[3] ), .d(\hdr_hld/low/U1664/U30/Z ), .e(
        \hdr_hld/low/U1664/x[2] ), .f(\hdr_hld/low/U1664/U30/Z ) );
    inv_1 \hdr_hld/low/U1664/U30/U30/Uinv  ( .x(\hdr_hld/low/U1664/U30/Z ), 
        .a(\hdr_hld/low/U1664/y[1] ) );
    aoi222_1 \hdr_hld/low/U1664/U31/U30/U1  ( .x(\hdr_hld/low/U1664/x[1] ), 
        .a(\hdr_hld/low/ncd[3] ), .b(\hdr_hld/low/ncd[2] ), .c(
        \hdr_hld/low/ncd[3] ), .d(\hdr_hld/low/U1664/U31/Z ), .e(
        \hdr_hld/low/ncd[2] ), .f(\hdr_hld/low/U1664/U31/Z ) );
    inv_1 \hdr_hld/low/U1664/U31/U30/Uinv  ( .x(\hdr_hld/low/U1664/U31/Z ), 
        .a(\hdr_hld/low/U1664/x[1] ) );
    aoi222_1 \hdr_hld/low/U1664/U37/U30/U1  ( .x(\hdr_hld/low/localcd ), .a(
        \hdr_hld/low/U1664/y[0] ), .b(\hdr_hld/low/U1664/y[1] ), .c(
        \hdr_hld/low/U1664/y[0] ), .d(\hdr_hld/low/U1664/U37/Z ), .e(
        \hdr_hld/low/U1664/y[1] ), .f(\hdr_hld/low/U1664/U37/Z ) );
    inv_1 \hdr_hld/low/U1664/U37/U30/Uinv  ( .x(\hdr_hld/low/U1664/U37/Z ), 
        .a(\hdr_hld/low/localcd ) );
    nor3_1 \hdr_hld/low/U1669/Unr  ( .x(\hdr_hld/low/U1669/nr ), .a(
        \hdr_hld/low/ctrlack_internal ), .b(\hdr_hld/low/driveh ), .c(n1) );
    nand3_1 \hdr_hld/low/U1669/Und  ( .x(\hdr_hld/low/U1669/nd ), .a(
        \hdr_hld/low/ctrlack_internal ), .b(n2), .c(\hdr_hld/low/drivel ) );
    oa21_1 \hdr_hld/low/U1669/U1  ( .x(\hdr_hld/low/U1669/n2 ), .a(
        \hdr_hld/low/U1669/n2 ), .b(\hdr_hld/low/U1669/nr ), .c(
        \hdr_hld/low/U1669/nd ) );
    inv_2 \hdr_hld/low/U1669/U3  ( .x(addr_req), .a(\hdr_hld/low/U1669/n2 ) );
    buf_2 \hdr_hld/high/U1653  ( .x(\hdr_hld/high/latch ), .a(\hdr_hld/net33 )
         );
    nor2_1 \hdr_hld/high/U264/U5  ( .x(\hdr_hld/high/nlocalcd ), .a(reset), 
        .b(\hdr_hld/high/localcd ) );
    nor2_1 \hdr_hld/high/U1659_0_/U5  ( .x(\hdr_hld/high/ncd[0] ), .a(itag_l
        [0]), .b(itag_h[0]) );
    nor2_1 \hdr_hld/high/U1659_1_/U5  ( .x(\hdr_hld/high/ncd[1] ), .a(itag_l
        [1]), .b(itag_h[1]) );
    nor2_1 \hdr_hld/high/U1659_2_/U5  ( .x(\hdr_hld/high/ncd[2] ), .a(itag_l
        [2]), .b(itag_h[2]) );
    nor2_1 \hdr_hld/high/U1659_3_/U5  ( .x(\hdr_hld/high/ncd[3] ), .a(itag_l
        [3]), .b(itag_h[3]) );
    nor2_1 \hdr_hld/high/U1659_4_/U5  ( .x(\hdr_hld/high/ncd[4] ), .a(itag_l
        [4]), .b(itag_h[4]) );
    nor2_1 \hdr_hld/high/U1659_5_/U5  ( .x(\hdr_hld/high/ncd[5] ), .a(col_l[0]
        ), .b(col_h[0]) );
    nor2_1 \hdr_hld/high/U1659_6_/U5  ( .x(\hdr_hld/high/ncd[6] ), .a(col_l[1]
        ), .b(col_h[1]) );
    nor2_1 \hdr_hld/high/U1659_7_/U5  ( .x(\hdr_hld/high/ncd[7] ), .a(col_l[2]
        ), .b(col_h[2]) );
    nor2_1 \hdr_hld/high/U3/U5  ( .x(\hdr_hld/high/ctrlack_internal ), .a(
        \hdr_hld/high/acb ), .b(\hdr_hld/high/ba ) );
    buf_2 \hdr_hld/high/U1665/U7  ( .x(\hdr_hld/high/driveh ), .a(receive) );
    buf_2 \hdr_hld/high/U1666/U7  ( .x(\hdr_hld/high/drivel ), .a(receive) );
    ao23_1 \hdr_hld/high/U1658_0_/U21/U1/U1  ( .x(itag_l[0]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[0]), .c(\hdr_hld/high/drivel ), .d(
        chwl[0]), .e(n7) );
    ao23_1 \hdr_hld/high/U1658_1_/U21/U1/U1  ( .x(itag_l[1]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[1]), .c(\hdr_hld/high/drivel ), .d(
        chwl[1]), .e(n7) );
    ao23_1 \hdr_hld/high/U1658_2_/U21/U1/U1  ( .x(itag_l[2]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[2]), .c(\hdr_hld/high/drivel ), .d(
        chwl[2]), .e(n7) );
    ao23_1 \hdr_hld/high/U1658_3_/U21/U1/U1  ( .x(itag_l[3]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[3]), .c(\hdr_hld/high/drivel ), .d(
        chwl[3]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1658_4_/U21/U1/U1  ( .x(itag_l[4]), .a(n4), .b(
        itag_l[4]), .c(\hdr_hld/high/drivel ), .d(chwl[4]), .e(
        \hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1658_5_/U21/U1/U1  ( .x(col_l[0]), .a(n4), .b(col_l
        [0]), .c(\hdr_hld/high/drivel ), .d(chwl[5]), .e(\hdr_hld/high/latch )
         );
    ao23_1 \hdr_hld/high/U1658_6_/U21/U1/U1  ( .x(col_l[1]), .a(
        \hdr_hld/high/drivel ), .b(col_l[1]), .c(\hdr_hld/high/drivel ), .d(
        chwl[6]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1658_7_/U21/U1/U1  ( .x(col_l[2]), .a(n4), .b(col_l
        [2]), .c(\hdr_hld/high/drivel ), .d(chwl[7]), .e(\hdr_hld/high/latch )
         );
    ao23_1 \hdr_hld/high/U1651_0_/U21/U1/U1  ( .x(itag_h[0]), .a(n5), .b(
        itag_h[0]), .c(n5), .d(chwh[0]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_1_/U21/U1/U1  ( .x(itag_h[1]), .a(n5), .b(
        itag_h[1]), .c(n6), .d(chwh[1]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_2_/U21/U1/U1  ( .x(itag_h[2]), .a(n5), .b(
        itag_h[2]), .c(n6), .d(chwh[2]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_3_/U21/U1/U1  ( .x(itag_h[3]), .a(n5), .b(
        itag_h[3]), .c(n6), .d(chwh[3]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_4_/U21/U1/U1  ( .x(itag_h[4]), .a(n5), .b(
        itag_h[4]), .c(n6), .d(chwh[4]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_5_/U21/U1/U1  ( .x(col_h[0]), .a(n5), .b(col_h
        [0]), .c(n6), .d(chwh[5]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_6_/U21/U1/U1  ( .x(col_h[1]), .a(n5), .b(col_h
        [1]), .c(n5), .d(chwh[6]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_7_/U21/U1/U1  ( .x(col_h[2]), .a(n5), .b(col_h
        [2]), .c(n5), .d(chwh[7]), .e(\hdr_hld/high/latch ) );
    aoai211_1 \hdr_hld/high/U4/U28/U1/U1  ( .x(\hdr_hld/high/U4/U28/U1/clr ), 
        .a(receive), .b(\hdr_hld/high/acb ), .c(\hdr_hld/high/nlocalcd ), .d(
        \hdr_hld/net33 ) );
    nand3_1 \hdr_hld/high/U4/U28/U1/U2  ( .x(\hdr_hld/high/U4/U28/U1/set ), 
        .a(\hdr_hld/high/nlocalcd ), .b(receive), .c(\hdr_hld/high/acb ) );
    nand2_2 \hdr_hld/high/U4/U28/U1/U3  ( .x(\hdr_hld/net33 ), .a(
        \hdr_hld/high/U4/U28/U1/clr ), .b(\hdr_hld/high/U4/U28/U1/set ) );
    oai21_1 \hdr_hld/high/U1/U30/U1/U1  ( .x(\hdr_hld/high/acb ), .a(
        \hdr_hld/high/U1/Z ), .b(\hdr_hld/high/ba ), .c(receive) );
    inv_1 \hdr_hld/high/U1/U30/U1/U2  ( .x(\hdr_hld/high/U1/Z ), .a(
        \hdr_hld/high/acb ) );
    ao222_1 \hdr_hld/high/U5/U18/U1/U1  ( .x(\hdr_hld/high/ba ), .a(
        \hdr_hld/high/latch ), .b(n9), .c(\hdr_hld/high/latch ), .d(
        \hdr_hld/high/ba ), .e(n9), .f(\hdr_hld/high/ba ) );
    aoi222_1 \hdr_hld/high/U1664/U28/U30/U1  ( .x(\hdr_hld/high/U1664/x[3] ), 
        .a(\hdr_hld/high/ncd[7] ), .b(\hdr_hld/high/ncd[6] ), .c(
        \hdr_hld/high/ncd[7] ), .d(\hdr_hld/high/U1664/U28/Z ), .e(
        \hdr_hld/high/ncd[6] ), .f(\hdr_hld/high/U1664/U28/Z ) );
    inv_1 \hdr_hld/high/U1664/U28/U30/Uinv  ( .x(\hdr_hld/high/U1664/U28/Z ), 
        .a(\hdr_hld/high/U1664/x[3] ) );
    aoi222_1 \hdr_hld/high/U1664/U32/U30/U1  ( .x(\hdr_hld/high/U1664/x[0] ), 
        .a(\hdr_hld/high/ncd[1] ), .b(\hdr_hld/high/ncd[0] ), .c(
        \hdr_hld/high/ncd[1] ), .d(\hdr_hld/high/U1664/U32/Z ), .e(
        \hdr_hld/high/ncd[0] ), .f(\hdr_hld/high/U1664/U32/Z ) );
    inv_1 \hdr_hld/high/U1664/U32/U30/Uinv  ( .x(\hdr_hld/high/U1664/U32/Z ), 
        .a(\hdr_hld/high/U1664/x[0] ) );
    aoi222_1 \hdr_hld/high/U1664/U29/U30/U1  ( .x(\hdr_hld/high/U1664/x[2] ), 
        .a(\hdr_hld/high/ncd[5] ), .b(\hdr_hld/high/ncd[4] ), .c(
        \hdr_hld/high/ncd[5] ), .d(\hdr_hld/high/U1664/U29/Z ), .e(
        \hdr_hld/high/ncd[4] ), .f(\hdr_hld/high/U1664/U29/Z ) );
    inv_1 \hdr_hld/high/U1664/U29/U30/Uinv  ( .x(\hdr_hld/high/U1664/U29/Z ), 
        .a(\hdr_hld/high/U1664/x[2] ) );
    aoi222_1 \hdr_hld/high/U1664/U33/U30/U1  ( .x(\hdr_hld/high/U1664/y[0] ), 
        .a(\hdr_hld/high/U1664/x[1] ), .b(\hdr_hld/high/U1664/x[0] ), .c(
        \hdr_hld/high/U1664/x[1] ), .d(\hdr_hld/high/U1664/U33/Z ), .e(
        \hdr_hld/high/U1664/x[0] ), .f(\hdr_hld/high/U1664/U33/Z ) );
    inv_1 \hdr_hld/high/U1664/U33/U30/Uinv  ( .x(\hdr_hld/high/U1664/U33/Z ), 
        .a(\hdr_hld/high/U1664/y[0] ) );
    aoi222_1 \hdr_hld/high/U1664/U30/U30/U1  ( .x(\hdr_hld/high/U1664/y[1] ), 
        .a(\hdr_hld/high/U1664/x[3] ), .b(\hdr_hld/high/U1664/x[2] ), .c(
        \hdr_hld/high/U1664/x[3] ), .d(\hdr_hld/high/U1664/U30/Z ), .e(
        \hdr_hld/high/U1664/x[2] ), .f(\hdr_hld/high/U1664/U30/Z ) );
    inv_1 \hdr_hld/high/U1664/U30/U30/Uinv  ( .x(\hdr_hld/high/U1664/U30/Z ), 
        .a(\hdr_hld/high/U1664/y[1] ) );
    aoi222_1 \hdr_hld/high/U1664/U31/U30/U1  ( .x(\hdr_hld/high/U1664/x[1] ), 
        .a(\hdr_hld/high/ncd[3] ), .b(\hdr_hld/high/ncd[2] ), .c(
        \hdr_hld/high/ncd[3] ), .d(\hdr_hld/high/U1664/U31/Z ), .e(
        \hdr_hld/high/ncd[2] ), .f(\hdr_hld/high/U1664/U31/Z ) );
    inv_1 \hdr_hld/high/U1664/U31/U30/Uinv  ( .x(\hdr_hld/high/U1664/U31/Z ), 
        .a(\hdr_hld/high/U1664/x[1] ) );
    aoi222_1 \hdr_hld/high/U1664/U37/U30/U1  ( .x(\hdr_hld/high/localcd ), .a(
        \hdr_hld/high/U1664/y[0] ), .b(\hdr_hld/high/U1664/y[1] ), .c(
        \hdr_hld/high/U1664/y[0] ), .d(\hdr_hld/high/U1664/U37/Z ), .e(
        \hdr_hld/high/U1664/y[1] ), .f(\hdr_hld/high/U1664/U37/Z ) );
    inv_1 \hdr_hld/high/U1664/U37/U30/Uinv  ( .x(\hdr_hld/high/U1664/U37/Z ), 
        .a(\hdr_hld/high/localcd ) );
    nor3_1 \hdr_hld/high/U1669/Unr  ( .x(\hdr_hld/high/U1669/nr ), .a(
        \hdr_hld/high/ctrlack_internal ), .b(\hdr_hld/high/drivel ), .c(n6) );
    nand3_1 \hdr_hld/high/U1669/Und  ( .x(\hdr_hld/high/U1669/nd ), .a(
        \hdr_hld/high/ctrlack_internal ), .b(\hdr_hld/high/drivel ), .c(n6) );
    oa21_1 \hdr_hld/high/U1669/U1  ( .x(\hdr_hld/high/U1669/n2 ), .a(
        \hdr_hld/high/U1669/n2 ), .b(\hdr_hld/high/U1669/nr ), .c(
        \hdr_hld/high/U1669/nd ) );
    inv_2 \hdr_hld/high/U1669/U3  ( .x(\hdr_hld/net20 ), .a(
        \hdr_hld/high/U1669/n2 ) );
    buf_2 U1 ( .x(n2), .a(\hdr_hld/net20 ) );
    buf_2 U2 ( .x(n1), .a(\hdr_hld/net20 ) );
    buf_1 U3 ( .x(n3), .a(\hdr_hld/low/latch ) );
    buf_1 U4 ( .x(n4), .a(\hdr_hld/high/drivel ) );
    buf_3 U5 ( .x(n5), .a(\hdr_hld/high/driveh ) );
    buf_3 U6 ( .x(n6), .a(\hdr_hld/high/driveh ) );
    buf_1 U7 ( .x(n7), .a(\hdr_hld/high/latch ) );
    inv_2 U8 ( .x(reset), .a(nReset) );
    buf_3 U9 ( .x(pullcd), .a(n9) );
endmodule


module chain_irdemux_32new_2 ( ctrlack, oh, ol, pullreq, pull_h, pull_l, 
    pullcd, reset, ctrlreq );
output [31:0] oh;
output [31:0] ol;
input  [7:0] pull_h;
input  [7:0] pull_l;
input  pullcd, reset, ctrlreq;
output ctrlack, pullreq;
    wire net30, net31, net17, \I0/net20 , \I0/net33 , \I0/net32 , 
        \I0/low/drivel , \I0/low/driveh , \I0/low/localcd , \I0/low/ncd[7] , 
        \I0/low/ncd[6] , \I0/low/ncd[5] , \I0/low/ncd[4] , \I0/low/ncd[3] , 
        \I0/low/ncd[2] , \I0/low/ncd[1] , \I0/low/ncd[0] , \I0/low/ba , 
        \I0/low/latch , \I0/low/acb , \I0/low/ctrlack_internal , 
        \I0/low/nlocalcd , \I0/low/U4/U28/U1/clr , \I0/low/U4/U28/U1/set , 
        \I0/low/U1/Z , \I0/low/U1664/y[0] , \I0/low/U1664/y[1] , 
        \I0/low/U1664/x[1] , \I0/low/U1664/x[3] , \I0/low/U1664/x[2] , 
        \I0/low/U1664/x[0] , \I0/low/U1664/U28/Z , \I0/low/U1664/U32/Z , 
        \I0/low/U1664/U29/Z , \I0/low/U1664/U33/Z , \I0/low/U1664/U30/Z , 
        \I0/low/U1664/U31/Z , \I0/low/U1664/U37/Z , \I0/low/U1669/nr , 
        \I0/low/U1669/nd , \I0/low/U1669/n2 , \I0/high/drivel , 
        \I0/high/driveh , \I0/high/localcd , \I0/high/ncd[7] , 
        \I0/high/ncd[6] , \I0/high/ncd[5] , \I0/high/ncd[4] , \I0/high/ncd[3] , 
        \I0/high/ncd[2] , \I0/high/ncd[1] , \I0/high/ncd[0] , \I0/high/ba , 
        \I0/high/latch , \I0/high/acb , \I0/high/ctrlack_internal , 
        \I0/high/nlocalcd , \I0/high/U4/U28/U1/clr , \I0/high/U4/U28/U1/set , 
        \I0/high/U1/Z , \I0/high/U1664/y[0] , \I0/high/U1664/y[1] , 
        \I0/high/U1664/x[1] , \I0/high/U1664/x[3] , \I0/high/U1664/x[2] , 
        \I0/high/U1664/x[0] , \I0/high/U1664/U28/Z , \I0/high/U1664/U32/Z , 
        \I0/high/U1664/U29/Z , \I0/high/U1664/U33/Z , \I0/high/U1664/U30/Z , 
        \I0/high/U1664/U31/Z , \I0/high/U1664/U37/Z , \I0/high/U1669/nr , 
        \I0/high/U1669/nd , \I0/high/U1669/n2 , \I1/net20 , \I1/net33 , 
        \I1/net32 , \I1/low/drivel , \I1/low/driveh , \I1/low/localcd , 
        \I1/low/ncd[7] , \I1/low/ncd[6] , \I1/low/ncd[5] , \I1/low/ncd[4] , 
        \I1/low/ncd[3] , \I1/low/ncd[2] , \I1/low/ncd[1] , \I1/low/ncd[0] , 
        \I1/low/ba , \I1/low/latch , \I1/low/acb , \I1/low/ctrlack_internal , 
        \I1/low/nlocalcd , \I1/low/U4/U28/U1/clr , \I1/low/U4/U28/U1/set , 
        \I1/low/U1/Z , \I1/low/U1664/y[0] , \I1/low/U1664/y[1] , 
        \I1/low/U1664/x[1] , \I1/low/U1664/x[3] , \I1/low/U1664/x[2] , 
        \I1/low/U1664/x[0] , \I1/low/U1664/U28/Z , \I1/low/U1664/U32/Z , 
        \I1/low/U1664/U29/Z , \I1/low/U1664/U33/Z , \I1/low/U1664/U30/Z , 
        \I1/low/U1664/U31/Z , \I1/low/U1664/U37/Z , \I1/low/U1669/nr , 
        \I1/low/U1669/nd , \I1/low/U1669/n2 , \I1/high/drivel , 
        \I1/high/driveh , \I1/high/localcd , \I1/high/ncd[7] , 
        \I1/high/ncd[6] , \I1/high/ncd[5] , \I1/high/ncd[4] , \I1/high/ncd[3] , 
        \I1/high/ncd[2] , \I1/high/ncd[1] , \I1/high/ncd[0] , \I1/high/ba , 
        \I1/high/latch , \I1/high/acb , \I1/high/ctrlack_internal , 
        \I1/high/nlocalcd , \I1/high/U4/U28/U1/clr , \I1/high/U4/U28/U1/set , 
        \I1/high/U1/Z , \I1/high/U1664/y[0] , \I1/high/U1664/y[1] , 
        \I1/high/U1664/x[1] , \I1/high/U1664/x[3] , \I1/high/U1664/x[2] , 
        \I1/high/U1664/x[0] , \I1/high/U1664/U28/Z , \I1/high/U1664/U32/Z , 
        \I1/high/U1664/U29/Z , \I1/high/U1664/U33/Z , \I1/high/U1664/U30/Z , 
        \I1/high/U1664/U31/Z , \I1/high/U1664/U37/Z , \I1/high/U1669/nr , 
        \I1/high/U1669/nd , \I1/high/U1669/n2 , n1, n2, n3, n4, n5, n6, n7, n8;
    nand2_1 \U3/U5  ( .x(pullreq), .a(net30), .b(net31) );
    nor2_1 \I0/U3/U5  ( .x(net30), .a(\I0/net32 ), .b(\I0/net33 ) );
    buf_2 \I0/low/U1653  ( .x(\I0/low/latch ), .a(\I0/net32 ) );
    nor2_1 \I0/low/U264/U5  ( .x(\I0/low/nlocalcd ), .a(reset), .b(
        \I0/low/localcd ) );
    nor2_1 \I0/low/U1659_0_/U5  ( .x(\I0/low/ncd[0] ), .a(ol[0]), .b(oh[0]) );
    nor2_1 \I0/low/U1659_1_/U5  ( .x(\I0/low/ncd[1] ), .a(ol[1]), .b(oh[1]) );
    nor2_1 \I0/low/U1659_2_/U5  ( .x(\I0/low/ncd[2] ), .a(ol[2]), .b(oh[2]) );
    nor2_1 \I0/low/U1659_3_/U5  ( .x(\I0/low/ncd[3] ), .a(ol[3]), .b(oh[3]) );
    nor2_1 \I0/low/U1659_4_/U5  ( .x(\I0/low/ncd[4] ), .a(ol[4]), .b(oh[4]) );
    nor2_1 \I0/low/U1659_5_/U5  ( .x(\I0/low/ncd[5] ), .a(ol[5]), .b(oh[5]) );
    nor2_1 \I0/low/U1659_6_/U5  ( .x(\I0/low/ncd[6] ), .a(ol[6]), .b(oh[6]) );
    nor2_1 \I0/low/U1659_7_/U5  ( .x(\I0/low/ncd[7] ), .a(ol[7]), .b(oh[7]) );
    nor2_1 \I0/low/U3/U5  ( .x(\I0/low/ctrlack_internal ), .a(\I0/low/acb ), 
        .b(\I0/low/ba ) );
    buf_2 \I0/low/U1665/U7  ( .x(\I0/low/driveh ), .a(\I0/net20 ) );
    buf_2 \I0/low/U1666/U7  ( .x(\I0/low/drivel ), .a(\I0/net20 ) );
    ao23_1 \I0/low/U1658_0_/U21/U1/U1  ( .x(ol[0]), .a(\I0/low/driveh ), .b(ol
        [0]), .c(n1), .d(pull_l[0]), .e(n2) );
    ao23_1 \I0/low/U1658_1_/U21/U1/U1  ( .x(ol[1]), .a(\I0/low/drivel ), .b(ol
        [1]), .c(\I0/low/driveh ), .d(pull_l[1]), .e(n2) );
    ao23_1 \I0/low/U1658_2_/U21/U1/U1  ( .x(ol[2]), .a(\I0/low/drivel ), .b(ol
        [2]), .c(\I0/low/driveh ), .d(pull_l[2]), .e(n2) );
    ao23_1 \I0/low/U1658_3_/U21/U1/U1  ( .x(ol[3]), .a(\I0/low/driveh ), .b(ol
        [3]), .c(\I0/low/drivel ), .d(pull_l[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_4_/U21/U1/U1  ( .x(ol[4]), .a(n1), .b(ol[4]), .c(
        \I0/low/drivel ), .d(pull_l[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_5_/U21/U1/U1  ( .x(ol[5]), .a(\I0/low/driveh ), .b(ol
        [5]), .c(n1), .d(pull_l[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_6_/U21/U1/U1  ( .x(ol[6]), .a(\I0/low/drivel ), .b(ol
        [6]), .c(\I0/low/driveh ), .d(pull_l[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_7_/U21/U1/U1  ( .x(ol[7]), .a(n1), .b(ol[7]), .c(n1), 
        .d(pull_l[7]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_0_/U21/U1/U1  ( .x(oh[0]), .a(\I0/low/driveh ), .b(oh
        [0]), .c(n1), .d(pull_h[0]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_1_/U21/U1/U1  ( .x(oh[1]), .a(n1), .b(oh[1]), .c(
        \I0/low/drivel ), .d(pull_h[1]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_2_/U21/U1/U1  ( .x(oh[2]), .a(\I0/low/drivel ), .b(oh
        [2]), .c(\I0/low/drivel ), .d(pull_h[2]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_3_/U21/U1/U1  ( .x(oh[3]), .a(n1), .b(oh[3]), .c(
        \I0/low/driveh ), .d(pull_h[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_4_/U21/U1/U1  ( .x(oh[4]), .a(n1), .b(oh[4]), .c(n1), 
        .d(pull_h[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_5_/U21/U1/U1  ( .x(oh[5]), .a(\I0/low/drivel ), .b(oh
        [5]), .c(n1), .d(pull_h[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_6_/U21/U1/U1  ( .x(oh[6]), .a(\I0/low/drivel ), .b(oh
        [6]), .c(\I0/low/driveh ), .d(pull_h[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_7_/U21/U1/U1  ( .x(oh[7]), .a(\I0/low/driveh ), .b(oh
        [7]), .c(\I0/low/drivel ), .d(pull_h[7]), .e(\I0/low/latch ) );
    aoai211_1 \I0/low/U4/U28/U1/U1  ( .x(\I0/low/U4/U28/U1/clr ), .a(
        \I0/net20 ), .b(\I0/low/acb ), .c(\I0/low/nlocalcd ), .d(\I0/net32 )
         );
    nand3_1 \I0/low/U4/U28/U1/U2  ( .x(\I0/low/U4/U28/U1/set ), .a(
        \I0/low/nlocalcd ), .b(\I0/net20 ), .c(\I0/low/acb ) );
    nand2_2 \I0/low/U4/U28/U1/U3  ( .x(\I0/net32 ), .a(\I0/low/U4/U28/U1/clr ), 
        .b(\I0/low/U4/U28/U1/set ) );
    oai21_1 \I0/low/U1/U30/U1/U1  ( .x(\I0/low/acb ), .a(\I0/low/U1/Z ), .b(
        \I0/low/ba ), .c(\I0/net20 ) );
    inv_1 \I0/low/U1/U30/U1/U2  ( .x(\I0/low/U1/Z ), .a(\I0/low/acb ) );
    ao222_1 \I0/low/U5/U18/U1/U1  ( .x(\I0/low/ba ), .a(\I0/low/latch ), .b(
        pullcd), .c(\I0/low/latch ), .d(\I0/low/ba ), .e(pullcd), .f(
        \I0/low/ba ) );
    aoi222_1 \I0/low/U1664/U28/U30/U1  ( .x(\I0/low/U1664/x[3] ), .a(
        \I0/low/ncd[7] ), .b(\I0/low/ncd[6] ), .c(\I0/low/ncd[7] ), .d(
        \I0/low/U1664/U28/Z ), .e(\I0/low/ncd[6] ), .f(\I0/low/U1664/U28/Z )
         );
    inv_1 \I0/low/U1664/U28/U30/Uinv  ( .x(\I0/low/U1664/U28/Z ), .a(
        \I0/low/U1664/x[3] ) );
    aoi222_1 \I0/low/U1664/U32/U30/U1  ( .x(\I0/low/U1664/x[0] ), .a(
        \I0/low/ncd[1] ), .b(\I0/low/ncd[0] ), .c(\I0/low/ncd[1] ), .d(
        \I0/low/U1664/U32/Z ), .e(\I0/low/ncd[0] ), .f(\I0/low/U1664/U32/Z )
         );
    inv_1 \I0/low/U1664/U32/U30/Uinv  ( .x(\I0/low/U1664/U32/Z ), .a(
        \I0/low/U1664/x[0] ) );
    aoi222_1 \I0/low/U1664/U29/U30/U1  ( .x(\I0/low/U1664/x[2] ), .a(
        \I0/low/ncd[5] ), .b(\I0/low/ncd[4] ), .c(\I0/low/ncd[5] ), .d(
        \I0/low/U1664/U29/Z ), .e(\I0/low/ncd[4] ), .f(\I0/low/U1664/U29/Z )
         );
    inv_1 \I0/low/U1664/U29/U30/Uinv  ( .x(\I0/low/U1664/U29/Z ), .a(
        \I0/low/U1664/x[2] ) );
    aoi222_1 \I0/low/U1664/U33/U30/U1  ( .x(\I0/low/U1664/y[0] ), .a(
        \I0/low/U1664/x[1] ), .b(\I0/low/U1664/x[0] ), .c(\I0/low/U1664/x[1] ), 
        .d(\I0/low/U1664/U33/Z ), .e(\I0/low/U1664/x[0] ), .f(
        \I0/low/U1664/U33/Z ) );
    inv_1 \I0/low/U1664/U33/U30/Uinv  ( .x(\I0/low/U1664/U33/Z ), .a(
        \I0/low/U1664/y[0] ) );
    aoi222_1 \I0/low/U1664/U30/U30/U1  ( .x(\I0/low/U1664/y[1] ), .a(
        \I0/low/U1664/x[3] ), .b(\I0/low/U1664/x[2] ), .c(\I0/low/U1664/x[3] ), 
        .d(\I0/low/U1664/U30/Z ), .e(\I0/low/U1664/x[2] ), .f(
        \I0/low/U1664/U30/Z ) );
    inv_1 \I0/low/U1664/U30/U30/Uinv  ( .x(\I0/low/U1664/U30/Z ), .a(
        \I0/low/U1664/y[1] ) );
    aoi222_1 \I0/low/U1664/U31/U30/U1  ( .x(\I0/low/U1664/x[1] ), .a(
        \I0/low/ncd[3] ), .b(\I0/low/ncd[2] ), .c(\I0/low/ncd[3] ), .d(
        \I0/low/U1664/U31/Z ), .e(\I0/low/ncd[2] ), .f(\I0/low/U1664/U31/Z )
         );
    inv_1 \I0/low/U1664/U31/U30/Uinv  ( .x(\I0/low/U1664/U31/Z ), .a(
        \I0/low/U1664/x[1] ) );
    aoi222_1 \I0/low/U1664/U37/U30/U1  ( .x(\I0/low/localcd ), .a(
        \I0/low/U1664/y[0] ), .b(\I0/low/U1664/y[1] ), .c(\I0/low/U1664/y[0] ), 
        .d(\I0/low/U1664/U37/Z ), .e(\I0/low/U1664/y[1] ), .f(
        \I0/low/U1664/U37/Z ) );
    inv_1 \I0/low/U1664/U37/U30/Uinv  ( .x(\I0/low/U1664/U37/Z ), .a(
        \I0/low/localcd ) );
    nor3_1 \I0/low/U1669/Unr  ( .x(\I0/low/U1669/nr ), .a(
        \I0/low/ctrlack_internal ), .b(n1), .c(\I0/low/driveh ) );
    nand3_1 \I0/low/U1669/Und  ( .x(\I0/low/U1669/nd ), .a(
        \I0/low/ctrlack_internal ), .b(\I0/low/drivel ), .c(\I0/low/driveh )
         );
    oa21_1 \I0/low/U1669/U1  ( .x(\I0/low/U1669/n2 ), .a(\I0/low/U1669/n2 ), 
        .b(\I0/low/U1669/nr ), .c(\I0/low/U1669/nd ) );
    inv_2 \I0/low/U1669/U3  ( .x(ctrlack), .a(\I0/low/U1669/n2 ) );
    buf_2 \I0/high/U1653  ( .x(\I0/high/latch ), .a(\I0/net33 ) );
    nor2_1 \I0/high/U264/U5  ( .x(\I0/high/nlocalcd ), .a(reset), .b(
        \I0/high/localcd ) );
    nor2_1 \I0/high/U1659_0_/U5  ( .x(\I0/high/ncd[0] ), .a(ol[8]), .b(oh[8])
         );
    nor2_1 \I0/high/U1659_1_/U5  ( .x(\I0/high/ncd[1] ), .a(ol[9]), .b(oh[9])
         );
    nor2_1 \I0/high/U1659_2_/U5  ( .x(\I0/high/ncd[2] ), .a(ol[10]), .b(oh[10]
        ) );
    nor2_1 \I0/high/U1659_3_/U5  ( .x(\I0/high/ncd[3] ), .a(ol[11]), .b(oh[11]
        ) );
    nor2_1 \I0/high/U1659_4_/U5  ( .x(\I0/high/ncd[4] ), .a(ol[12]), .b(oh[12]
        ) );
    nor2_1 \I0/high/U1659_5_/U5  ( .x(\I0/high/ncd[5] ), .a(ol[13]), .b(oh[13]
        ) );
    nor2_1 \I0/high/U1659_6_/U5  ( .x(\I0/high/ncd[6] ), .a(ol[14]), .b(oh[14]
        ) );
    nor2_1 \I0/high/U1659_7_/U5  ( .x(\I0/high/ncd[7] ), .a(ol[15]), .b(oh[15]
        ) );
    nor2_1 \I0/high/U3/U5  ( .x(\I0/high/ctrlack_internal ), .a(\I0/high/acb ), 
        .b(\I0/high/ba ) );
    buf_2 \I0/high/U1665/U7  ( .x(\I0/high/driveh ), .a(net17) );
    buf_2 \I0/high/U1666/U7  ( .x(\I0/high/drivel ), .a(net17) );
    ao23_1 \I0/high/U1658_0_/U21/U1/U1  ( .x(ol[8]), .a(\I0/high/driveh ), .b(
        ol[8]), .c(n3), .d(pull_l[0]), .e(n4) );
    ao23_1 \I0/high/U1658_1_/U21/U1/U1  ( .x(ol[9]), .a(\I0/high/drivel ), .b(
        ol[9]), .c(\I0/high/driveh ), .d(pull_l[1]), .e(n4) );
    ao23_1 \I0/high/U1658_2_/U21/U1/U1  ( .x(ol[10]), .a(\I0/high/drivel ), 
        .b(ol[10]), .c(\I0/high/driveh ), .d(pull_l[2]), .e(n4) );
    ao23_1 \I0/high/U1658_3_/U21/U1/U1  ( .x(ol[11]), .a(\I0/high/driveh ), 
        .b(ol[11]), .c(\I0/high/drivel ), .d(pull_l[3]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_4_/U21/U1/U1  ( .x(ol[12]), .a(n3), .b(ol[12]), .c(
        \I0/high/drivel ), .d(pull_l[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_5_/U21/U1/U1  ( .x(ol[13]), .a(\I0/high/driveh ), 
        .b(ol[13]), .c(n3), .d(pull_l[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_6_/U21/U1/U1  ( .x(ol[14]), .a(\I0/high/drivel ), 
        .b(ol[14]), .c(\I0/high/driveh ), .d(pull_l[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_7_/U21/U1/U1  ( .x(ol[15]), .a(n3), .b(ol[15]), .c(
        n3), .d(pull_l[7]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_0_/U21/U1/U1  ( .x(oh[8]), .a(\I0/high/driveh ), .b(
        oh[8]), .c(n3), .d(pull_h[0]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_1_/U21/U1/U1  ( .x(oh[9]), .a(n3), .b(oh[9]), .c(
        \I0/high/drivel ), .d(pull_h[1]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_2_/U21/U1/U1  ( .x(oh[10]), .a(\I0/high/drivel ), 
        .b(oh[10]), .c(\I0/high/drivel ), .d(pull_h[2]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_3_/U21/U1/U1  ( .x(oh[11]), .a(n3), .b(oh[11]), .c(
        \I0/high/driveh ), .d(pull_h[3]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_4_/U21/U1/U1  ( .x(oh[12]), .a(n3), .b(oh[12]), .c(
        n3), .d(pull_h[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_5_/U21/U1/U1  ( .x(oh[13]), .a(\I0/high/drivel ), 
        .b(oh[13]), .c(n3), .d(pull_h[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_6_/U21/U1/U1  ( .x(oh[14]), .a(\I0/high/drivel ), 
        .b(oh[14]), .c(\I0/high/driveh ), .d(pull_h[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_7_/U21/U1/U1  ( .x(oh[15]), .a(\I0/high/driveh ), 
        .b(oh[15]), .c(\I0/high/drivel ), .d(pull_h[7]), .e(\I0/high/latch )
         );
    aoai211_1 \I0/high/U4/U28/U1/U1  ( .x(\I0/high/U4/U28/U1/clr ), .a(net17), 
        .b(\I0/high/acb ), .c(\I0/high/nlocalcd ), .d(\I0/net33 ) );
    nand3_1 \I0/high/U4/U28/U1/U2  ( .x(\I0/high/U4/U28/U1/set ), .a(
        \I0/high/nlocalcd ), .b(net17), .c(\I0/high/acb ) );
    nand2_2 \I0/high/U4/U28/U1/U3  ( .x(\I0/net33 ), .a(
        \I0/high/U4/U28/U1/clr ), .b(\I0/high/U4/U28/U1/set ) );
    oai21_1 \I0/high/U1/U30/U1/U1  ( .x(\I0/high/acb ), .a(\I0/high/U1/Z ), 
        .b(\I0/high/ba ), .c(net17) );
    inv_1 \I0/high/U1/U30/U1/U2  ( .x(\I0/high/U1/Z ), .a(\I0/high/acb ) );
    ao222_1 \I0/high/U5/U18/U1/U1  ( .x(\I0/high/ba ), .a(\I0/high/latch ), 
        .b(pullcd), .c(\I0/high/latch ), .d(\I0/high/ba ), .e(pullcd), .f(
        \I0/high/ba ) );
    aoi222_1 \I0/high/U1664/U28/U30/U1  ( .x(\I0/high/U1664/x[3] ), .a(
        \I0/high/ncd[7] ), .b(\I0/high/ncd[6] ), .c(\I0/high/ncd[7] ), .d(
        \I0/high/U1664/U28/Z ), .e(\I0/high/ncd[6] ), .f(\I0/high/U1664/U28/Z 
        ) );
    inv_1 \I0/high/U1664/U28/U30/Uinv  ( .x(\I0/high/U1664/U28/Z ), .a(
        \I0/high/U1664/x[3] ) );
    aoi222_1 \I0/high/U1664/U32/U30/U1  ( .x(\I0/high/U1664/x[0] ), .a(
        \I0/high/ncd[1] ), .b(\I0/high/ncd[0] ), .c(\I0/high/ncd[1] ), .d(
        \I0/high/U1664/U32/Z ), .e(\I0/high/ncd[0] ), .f(\I0/high/U1664/U32/Z 
        ) );
    inv_1 \I0/high/U1664/U32/U30/Uinv  ( .x(\I0/high/U1664/U32/Z ), .a(
        \I0/high/U1664/x[0] ) );
    aoi222_1 \I0/high/U1664/U29/U30/U1  ( .x(\I0/high/U1664/x[2] ), .a(
        \I0/high/ncd[5] ), .b(\I0/high/ncd[4] ), .c(\I0/high/ncd[5] ), .d(
        \I0/high/U1664/U29/Z ), .e(\I0/high/ncd[4] ), .f(\I0/high/U1664/U29/Z 
        ) );
    inv_1 \I0/high/U1664/U29/U30/Uinv  ( .x(\I0/high/U1664/U29/Z ), .a(
        \I0/high/U1664/x[2] ) );
    aoi222_1 \I0/high/U1664/U33/U30/U1  ( .x(\I0/high/U1664/y[0] ), .a(
        \I0/high/U1664/x[1] ), .b(\I0/high/U1664/x[0] ), .c(
        \I0/high/U1664/x[1] ), .d(\I0/high/U1664/U33/Z ), .e(
        \I0/high/U1664/x[0] ), .f(\I0/high/U1664/U33/Z ) );
    inv_1 \I0/high/U1664/U33/U30/Uinv  ( .x(\I0/high/U1664/U33/Z ), .a(
        \I0/high/U1664/y[0] ) );
    aoi222_1 \I0/high/U1664/U30/U30/U1  ( .x(\I0/high/U1664/y[1] ), .a(
        \I0/high/U1664/x[3] ), .b(\I0/high/U1664/x[2] ), .c(
        \I0/high/U1664/x[3] ), .d(\I0/high/U1664/U30/Z ), .e(
        \I0/high/U1664/x[2] ), .f(\I0/high/U1664/U30/Z ) );
    inv_1 \I0/high/U1664/U30/U30/Uinv  ( .x(\I0/high/U1664/U30/Z ), .a(
        \I0/high/U1664/y[1] ) );
    aoi222_1 \I0/high/U1664/U31/U30/U1  ( .x(\I0/high/U1664/x[1] ), .a(
        \I0/high/ncd[3] ), .b(\I0/high/ncd[2] ), .c(\I0/high/ncd[3] ), .d(
        \I0/high/U1664/U31/Z ), .e(\I0/high/ncd[2] ), .f(\I0/high/U1664/U31/Z 
        ) );
    inv_1 \I0/high/U1664/U31/U30/Uinv  ( .x(\I0/high/U1664/U31/Z ), .a(
        \I0/high/U1664/x[1] ) );
    aoi222_1 \I0/high/U1664/U37/U30/U1  ( .x(\I0/high/localcd ), .a(
        \I0/high/U1664/y[0] ), .b(\I0/high/U1664/y[1] ), .c(
        \I0/high/U1664/y[0] ), .d(\I0/high/U1664/U37/Z ), .e(
        \I0/high/U1664/y[1] ), .f(\I0/high/U1664/U37/Z ) );
    inv_1 \I0/high/U1664/U37/U30/Uinv  ( .x(\I0/high/U1664/U37/Z ), .a(
        \I0/high/localcd ) );
    nor3_1 \I0/high/U1669/Unr  ( .x(\I0/high/U1669/nr ), .a(
        \I0/high/ctrlack_internal ), .b(n3), .c(\I0/high/driveh ) );
    nand3_1 \I0/high/U1669/Und  ( .x(\I0/high/U1669/nd ), .a(
        \I0/high/ctrlack_internal ), .b(\I0/high/drivel ), .c(\I0/high/driveh 
        ) );
    oa21_1 \I0/high/U1669/U1  ( .x(\I0/high/U1669/n2 ), .a(\I0/high/U1669/n2 ), 
        .b(\I0/high/U1669/nr ), .c(\I0/high/U1669/nd ) );
    inv_2 \I0/high/U1669/U3  ( .x(\I0/net20 ), .a(\I0/high/U1669/n2 ) );
    nor2_1 \I1/U3/U5  ( .x(net31), .a(\I1/net32 ), .b(\I1/net33 ) );
    buf_2 \I1/low/U1653  ( .x(\I1/low/latch ), .a(\I1/net32 ) );
    nor2_1 \I1/low/U264/U5  ( .x(\I1/low/nlocalcd ), .a(reset), .b(
        \I1/low/localcd ) );
    nor2_1 \I1/low/U1659_0_/U5  ( .x(\I1/low/ncd[0] ), .a(ol[16]), .b(oh[16])
         );
    nor2_1 \I1/low/U1659_1_/U5  ( .x(\I1/low/ncd[1] ), .a(ol[17]), .b(oh[17])
         );
    nor2_1 \I1/low/U1659_2_/U5  ( .x(\I1/low/ncd[2] ), .a(ol[18]), .b(oh[18])
         );
    nor2_1 \I1/low/U1659_3_/U5  ( .x(\I1/low/ncd[3] ), .a(ol[19]), .b(oh[19])
         );
    nor2_1 \I1/low/U1659_4_/U5  ( .x(\I1/low/ncd[4] ), .a(ol[20]), .b(oh[20])
         );
    nor2_1 \I1/low/U1659_5_/U5  ( .x(\I1/low/ncd[5] ), .a(ol[21]), .b(oh[21])
         );
    nor2_1 \I1/low/U1659_6_/U5  ( .x(\I1/low/ncd[6] ), .a(ol[22]), .b(oh[22])
         );
    nor2_1 \I1/low/U1659_7_/U5  ( .x(\I1/low/ncd[7] ), .a(ol[23]), .b(oh[23])
         );
    nor2_1 \I1/low/U3/U5  ( .x(\I1/low/ctrlack_internal ), .a(\I1/low/acb ), 
        .b(\I1/low/ba ) );
    buf_2 \I1/low/U1665/U7  ( .x(\I1/low/driveh ), .a(\I1/net20 ) );
    buf_2 \I1/low/U1666/U7  ( .x(\I1/low/drivel ), .a(\I1/net20 ) );
    ao23_1 \I1/low/U1658_0_/U21/U1/U1  ( .x(ol[16]), .a(\I1/low/driveh ), .b(
        ol[16]), .c(n5), .d(pull_l[0]), .e(n6) );
    ao23_1 \I1/low/U1658_1_/U21/U1/U1  ( .x(ol[17]), .a(\I1/low/drivel ), .b(
        ol[17]), .c(\I1/low/driveh ), .d(pull_l[1]), .e(n6) );
    ao23_1 \I1/low/U1658_2_/U21/U1/U1  ( .x(ol[18]), .a(\I1/low/drivel ), .b(
        ol[18]), .c(\I1/low/driveh ), .d(pull_l[2]), .e(n6) );
    ao23_1 \I1/low/U1658_3_/U21/U1/U1  ( .x(ol[19]), .a(\I1/low/driveh ), .b(
        ol[19]), .c(\I1/low/drivel ), .d(pull_l[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_4_/U21/U1/U1  ( .x(ol[20]), .a(n5), .b(ol[20]), .c(
        \I1/low/drivel ), .d(pull_l[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_5_/U21/U1/U1  ( .x(ol[21]), .a(\I1/low/driveh ), .b(
        ol[21]), .c(n5), .d(pull_l[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_6_/U21/U1/U1  ( .x(ol[22]), .a(\I1/low/drivel ), .b(
        ol[22]), .c(\I1/low/driveh ), .d(pull_l[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_7_/U21/U1/U1  ( .x(ol[23]), .a(n5), .b(ol[23]), .c(n5
        ), .d(pull_l[7]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_0_/U21/U1/U1  ( .x(oh[16]), .a(\I1/low/driveh ), .b(
        oh[16]), .c(n5), .d(pull_h[0]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_1_/U21/U1/U1  ( .x(oh[17]), .a(n5), .b(oh[17]), .c(
        \I1/low/drivel ), .d(pull_h[1]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_2_/U21/U1/U1  ( .x(oh[18]), .a(\I1/low/drivel ), .b(
        oh[18]), .c(\I1/low/drivel ), .d(pull_h[2]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_3_/U21/U1/U1  ( .x(oh[19]), .a(n5), .b(oh[19]), .c(
        \I1/low/driveh ), .d(pull_h[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_4_/U21/U1/U1  ( .x(oh[20]), .a(n5), .b(oh[20]), .c(n5
        ), .d(pull_h[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_5_/U21/U1/U1  ( .x(oh[21]), .a(\I1/low/drivel ), .b(
        oh[21]), .c(n5), .d(pull_h[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_6_/U21/U1/U1  ( .x(oh[22]), .a(\I1/low/drivel ), .b(
        oh[22]), .c(\I1/low/driveh ), .d(pull_h[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_7_/U21/U1/U1  ( .x(oh[23]), .a(\I1/low/driveh ), .b(
        oh[23]), .c(\I1/low/drivel ), .d(pull_h[7]), .e(\I1/low/latch ) );
    aoai211_1 \I1/low/U4/U28/U1/U1  ( .x(\I1/low/U4/U28/U1/clr ), .a(
        \I1/net20 ), .b(\I1/low/acb ), .c(\I1/low/nlocalcd ), .d(\I1/net32 )
         );
    nand3_1 \I1/low/U4/U28/U1/U2  ( .x(\I1/low/U4/U28/U1/set ), .a(
        \I1/low/nlocalcd ), .b(\I1/net20 ), .c(\I1/low/acb ) );
    nand2_2 \I1/low/U4/U28/U1/U3  ( .x(\I1/net32 ), .a(\I1/low/U4/U28/U1/clr ), 
        .b(\I1/low/U4/U28/U1/set ) );
    oai21_1 \I1/low/U1/U30/U1/U1  ( .x(\I1/low/acb ), .a(\I1/low/U1/Z ), .b(
        \I1/low/ba ), .c(\I1/net20 ) );
    inv_1 \I1/low/U1/U30/U1/U2  ( .x(\I1/low/U1/Z ), .a(\I1/low/acb ) );
    ao222_1 \I1/low/U5/U18/U1/U1  ( .x(\I1/low/ba ), .a(\I1/low/latch ), .b(
        pullcd), .c(\I1/low/latch ), .d(\I1/low/ba ), .e(pullcd), .f(
        \I1/low/ba ) );
    aoi222_1 \I1/low/U1664/U28/U30/U1  ( .x(\I1/low/U1664/x[3] ), .a(
        \I1/low/ncd[7] ), .b(\I1/low/ncd[6] ), .c(\I1/low/ncd[7] ), .d(
        \I1/low/U1664/U28/Z ), .e(\I1/low/ncd[6] ), .f(\I1/low/U1664/U28/Z )
         );
    inv_1 \I1/low/U1664/U28/U30/Uinv  ( .x(\I1/low/U1664/U28/Z ), .a(
        \I1/low/U1664/x[3] ) );
    aoi222_1 \I1/low/U1664/U32/U30/U1  ( .x(\I1/low/U1664/x[0] ), .a(
        \I1/low/ncd[1] ), .b(\I1/low/ncd[0] ), .c(\I1/low/ncd[1] ), .d(
        \I1/low/U1664/U32/Z ), .e(\I1/low/ncd[0] ), .f(\I1/low/U1664/U32/Z )
         );
    inv_1 \I1/low/U1664/U32/U30/Uinv  ( .x(\I1/low/U1664/U32/Z ), .a(
        \I1/low/U1664/x[0] ) );
    aoi222_1 \I1/low/U1664/U29/U30/U1  ( .x(\I1/low/U1664/x[2] ), .a(
        \I1/low/ncd[5] ), .b(\I1/low/ncd[4] ), .c(\I1/low/ncd[5] ), .d(
        \I1/low/U1664/U29/Z ), .e(\I1/low/ncd[4] ), .f(\I1/low/U1664/U29/Z )
         );
    inv_1 \I1/low/U1664/U29/U30/Uinv  ( .x(\I1/low/U1664/U29/Z ), .a(
        \I1/low/U1664/x[2] ) );
    aoi222_1 \I1/low/U1664/U33/U30/U1  ( .x(\I1/low/U1664/y[0] ), .a(
        \I1/low/U1664/x[1] ), .b(\I1/low/U1664/x[0] ), .c(\I1/low/U1664/x[1] ), 
        .d(\I1/low/U1664/U33/Z ), .e(\I1/low/U1664/x[0] ), .f(
        \I1/low/U1664/U33/Z ) );
    inv_1 \I1/low/U1664/U33/U30/Uinv  ( .x(\I1/low/U1664/U33/Z ), .a(
        \I1/low/U1664/y[0] ) );
    aoi222_1 \I1/low/U1664/U30/U30/U1  ( .x(\I1/low/U1664/y[1] ), .a(
        \I1/low/U1664/x[3] ), .b(\I1/low/U1664/x[2] ), .c(\I1/low/U1664/x[3] ), 
        .d(\I1/low/U1664/U30/Z ), .e(\I1/low/U1664/x[2] ), .f(
        \I1/low/U1664/U30/Z ) );
    inv_1 \I1/low/U1664/U30/U30/Uinv  ( .x(\I1/low/U1664/U30/Z ), .a(
        \I1/low/U1664/y[1] ) );
    aoi222_1 \I1/low/U1664/U31/U30/U1  ( .x(\I1/low/U1664/x[1] ), .a(
        \I1/low/ncd[3] ), .b(\I1/low/ncd[2] ), .c(\I1/low/ncd[3] ), .d(
        \I1/low/U1664/U31/Z ), .e(\I1/low/ncd[2] ), .f(\I1/low/U1664/U31/Z )
         );
    inv_1 \I1/low/U1664/U31/U30/Uinv  ( .x(\I1/low/U1664/U31/Z ), .a(
        \I1/low/U1664/x[1] ) );
    aoi222_1 \I1/low/U1664/U37/U30/U1  ( .x(\I1/low/localcd ), .a(
        \I1/low/U1664/y[0] ), .b(\I1/low/U1664/y[1] ), .c(\I1/low/U1664/y[0] ), 
        .d(\I1/low/U1664/U37/Z ), .e(\I1/low/U1664/y[1] ), .f(
        \I1/low/U1664/U37/Z ) );
    inv_1 \I1/low/U1664/U37/U30/Uinv  ( .x(\I1/low/U1664/U37/Z ), .a(
        \I1/low/localcd ) );
    nor3_1 \I1/low/U1669/Unr  ( .x(\I1/low/U1669/nr ), .a(
        \I1/low/ctrlack_internal ), .b(n5), .c(\I1/low/driveh ) );
    nand3_1 \I1/low/U1669/Und  ( .x(\I1/low/U1669/nd ), .a(
        \I1/low/ctrlack_internal ), .b(\I1/low/drivel ), .c(\I1/low/driveh )
         );
    oa21_1 \I1/low/U1669/U1  ( .x(\I1/low/U1669/n2 ), .a(\I1/low/U1669/n2 ), 
        .b(\I1/low/U1669/nr ), .c(\I1/low/U1669/nd ) );
    inv_2 \I1/low/U1669/U3  ( .x(net17), .a(\I1/low/U1669/n2 ) );
    buf_2 \I1/high/U1653  ( .x(\I1/high/latch ), .a(\I1/net33 ) );
    nor2_1 \I1/high/U264/U5  ( .x(\I1/high/nlocalcd ), .a(reset), .b(
        \I1/high/localcd ) );
    nor2_1 \I1/high/U1659_0_/U5  ( .x(\I1/high/ncd[0] ), .a(ol[24]), .b(oh[24]
        ) );
    nor2_1 \I1/high/U1659_1_/U5  ( .x(\I1/high/ncd[1] ), .a(ol[25]), .b(oh[25]
        ) );
    nor2_1 \I1/high/U1659_2_/U5  ( .x(\I1/high/ncd[2] ), .a(ol[26]), .b(oh[26]
        ) );
    nor2_1 \I1/high/U1659_3_/U5  ( .x(\I1/high/ncd[3] ), .a(ol[27]), .b(oh[27]
        ) );
    nor2_1 \I1/high/U1659_4_/U5  ( .x(\I1/high/ncd[4] ), .a(ol[28]), .b(oh[28]
        ) );
    nor2_1 \I1/high/U1659_5_/U5  ( .x(\I1/high/ncd[5] ), .a(ol[29]), .b(oh[29]
        ) );
    nor2_1 \I1/high/U1659_6_/U5  ( .x(\I1/high/ncd[6] ), .a(ol[30]), .b(oh[30]
        ) );
    nor2_1 \I1/high/U1659_7_/U5  ( .x(\I1/high/ncd[7] ), .a(ol[31]), .b(oh[31]
        ) );
    nor2_1 \I1/high/U3/U5  ( .x(\I1/high/ctrlack_internal ), .a(\I1/high/acb ), 
        .b(\I1/high/ba ) );
    buf_2 \I1/high/U1665/U7  ( .x(\I1/high/driveh ), .a(ctrlreq) );
    buf_2 \I1/high/U1666/U7  ( .x(\I1/high/drivel ), .a(ctrlreq) );
    ao23_1 \I1/high/U1658_0_/U21/U1/U1  ( .x(ol[24]), .a(\I1/high/driveh ), 
        .b(ol[24]), .c(n7), .d(pull_l[0]), .e(n8) );
    ao23_1 \I1/high/U1658_1_/U21/U1/U1  ( .x(ol[25]), .a(\I1/high/drivel ), 
        .b(ol[25]), .c(\I1/high/driveh ), .d(pull_l[1]), .e(n8) );
    ao23_1 \I1/high/U1658_2_/U21/U1/U1  ( .x(ol[26]), .a(\I1/high/drivel ), 
        .b(ol[26]), .c(\I1/high/driveh ), .d(pull_l[2]), .e(n8) );
    ao23_1 \I1/high/U1658_3_/U21/U1/U1  ( .x(ol[27]), .a(\I1/high/driveh ), 
        .b(ol[27]), .c(\I1/high/drivel ), .d(pull_l[3]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1658_4_/U21/U1/U1  ( .x(ol[28]), .a(n7), .b(ol[28]), .c(
        \I1/high/drivel ), .d(pull_l[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_5_/U21/U1/U1  ( .x(ol[29]), .a(\I1/high/driveh ), 
        .b(ol[29]), .c(n7), .d(pull_l[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_6_/U21/U1/U1  ( .x(ol[30]), .a(\I1/high/drivel ), 
        .b(ol[30]), .c(\I1/high/driveh ), .d(pull_l[6]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1658_7_/U21/U1/U1  ( .x(ol[31]), .a(n7), .b(ol[31]), .c(
        n7), .d(pull_l[7]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_0_/U21/U1/U1  ( .x(oh[24]), .a(\I1/high/driveh ), 
        .b(oh[24]), .c(n7), .d(pull_h[0]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_1_/U21/U1/U1  ( .x(oh[25]), .a(n7), .b(oh[25]), .c(
        \I1/high/drivel ), .d(pull_h[1]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_2_/U21/U1/U1  ( .x(oh[26]), .a(\I1/high/drivel ), 
        .b(oh[26]), .c(\I1/high/drivel ), .d(pull_h[2]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1651_3_/U21/U1/U1  ( .x(oh[27]), .a(n7), .b(oh[27]), .c(
        \I1/high/driveh ), .d(pull_h[3]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_4_/U21/U1/U1  ( .x(oh[28]), .a(n7), .b(oh[28]), .c(
        n7), .d(pull_h[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_5_/U21/U1/U1  ( .x(oh[29]), .a(\I1/high/drivel ), 
        .b(oh[29]), .c(n7), .d(pull_h[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_6_/U21/U1/U1  ( .x(oh[30]), .a(\I1/high/drivel ), 
        .b(oh[30]), .c(\I1/high/driveh ), .d(pull_h[6]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1651_7_/U21/U1/U1  ( .x(oh[31]), .a(\I1/high/driveh ), 
        .b(oh[31]), .c(\I1/high/drivel ), .d(pull_h[7]), .e(\I1/high/latch )
         );
    aoai211_1 \I1/high/U4/U28/U1/U1  ( .x(\I1/high/U4/U28/U1/clr ), .a(ctrlreq
        ), .b(\I1/high/acb ), .c(\I1/high/nlocalcd ), .d(\I1/net33 ) );
    nand3_1 \I1/high/U4/U28/U1/U2  ( .x(\I1/high/U4/U28/U1/set ), .a(
        \I1/high/nlocalcd ), .b(ctrlreq), .c(\I1/high/acb ) );
    nand2_2 \I1/high/U4/U28/U1/U3  ( .x(\I1/net33 ), .a(
        \I1/high/U4/U28/U1/clr ), .b(\I1/high/U4/U28/U1/set ) );
    oai21_1 \I1/high/U1/U30/U1/U1  ( .x(\I1/high/acb ), .a(\I1/high/U1/Z ), 
        .b(\I1/high/ba ), .c(ctrlreq) );
    inv_1 \I1/high/U1/U30/U1/U2  ( .x(\I1/high/U1/Z ), .a(\I1/high/acb ) );
    ao222_1 \I1/high/U5/U18/U1/U1  ( .x(\I1/high/ba ), .a(\I1/high/latch ), 
        .b(pullcd), .c(\I1/high/latch ), .d(\I1/high/ba ), .e(pullcd), .f(
        \I1/high/ba ) );
    aoi222_1 \I1/high/U1664/U28/U30/U1  ( .x(\I1/high/U1664/x[3] ), .a(
        \I1/high/ncd[7] ), .b(\I1/high/ncd[6] ), .c(\I1/high/ncd[7] ), .d(
        \I1/high/U1664/U28/Z ), .e(\I1/high/ncd[6] ), .f(\I1/high/U1664/U28/Z 
        ) );
    inv_1 \I1/high/U1664/U28/U30/Uinv  ( .x(\I1/high/U1664/U28/Z ), .a(
        \I1/high/U1664/x[3] ) );
    aoi222_1 \I1/high/U1664/U32/U30/U1  ( .x(\I1/high/U1664/x[0] ), .a(
        \I1/high/ncd[1] ), .b(\I1/high/ncd[0] ), .c(\I1/high/ncd[1] ), .d(
        \I1/high/U1664/U32/Z ), .e(\I1/high/ncd[0] ), .f(\I1/high/U1664/U32/Z 
        ) );
    inv_1 \I1/high/U1664/U32/U30/Uinv  ( .x(\I1/high/U1664/U32/Z ), .a(
        \I1/high/U1664/x[0] ) );
    aoi222_1 \I1/high/U1664/U29/U30/U1  ( .x(\I1/high/U1664/x[2] ), .a(
        \I1/high/ncd[5] ), .b(\I1/high/ncd[4] ), .c(\I1/high/ncd[5] ), .d(
        \I1/high/U1664/U29/Z ), .e(\I1/high/ncd[4] ), .f(\I1/high/U1664/U29/Z 
        ) );
    inv_1 \I1/high/U1664/U29/U30/Uinv  ( .x(\I1/high/U1664/U29/Z ), .a(
        \I1/high/U1664/x[2] ) );
    aoi222_1 \I1/high/U1664/U33/U30/U1  ( .x(\I1/high/U1664/y[0] ), .a(
        \I1/high/U1664/x[1] ), .b(\I1/high/U1664/x[0] ), .c(
        \I1/high/U1664/x[1] ), .d(\I1/high/U1664/U33/Z ), .e(
        \I1/high/U1664/x[0] ), .f(\I1/high/U1664/U33/Z ) );
    inv_1 \I1/high/U1664/U33/U30/Uinv  ( .x(\I1/high/U1664/U33/Z ), .a(
        \I1/high/U1664/y[0] ) );
    aoi222_1 \I1/high/U1664/U30/U30/U1  ( .x(\I1/high/U1664/y[1] ), .a(
        \I1/high/U1664/x[3] ), .b(\I1/high/U1664/x[2] ), .c(
        \I1/high/U1664/x[3] ), .d(\I1/high/U1664/U30/Z ), .e(
        \I1/high/U1664/x[2] ), .f(\I1/high/U1664/U30/Z ) );
    inv_1 \I1/high/U1664/U30/U30/Uinv  ( .x(\I1/high/U1664/U30/Z ), .a(
        \I1/high/U1664/y[1] ) );
    aoi222_1 \I1/high/U1664/U31/U30/U1  ( .x(\I1/high/U1664/x[1] ), .a(
        \I1/high/ncd[3] ), .b(\I1/high/ncd[2] ), .c(\I1/high/ncd[3] ), .d(
        \I1/high/U1664/U31/Z ), .e(\I1/high/ncd[2] ), .f(\I1/high/U1664/U31/Z 
        ) );
    inv_1 \I1/high/U1664/U31/U30/Uinv  ( .x(\I1/high/U1664/U31/Z ), .a(
        \I1/high/U1664/x[1] ) );
    aoi222_1 \I1/high/U1664/U37/U30/U1  ( .x(\I1/high/localcd ), .a(
        \I1/high/U1664/y[0] ), .b(\I1/high/U1664/y[1] ), .c(
        \I1/high/U1664/y[0] ), .d(\I1/high/U1664/U37/Z ), .e(
        \I1/high/U1664/y[1] ), .f(\I1/high/U1664/U37/Z ) );
    inv_1 \I1/high/U1664/U37/U30/Uinv  ( .x(\I1/high/U1664/U37/Z ), .a(
        \I1/high/localcd ) );
    nor3_1 \I1/high/U1669/Unr  ( .x(\I1/high/U1669/nr ), .a(
        \I1/high/ctrlack_internal ), .b(n7), .c(\I1/high/driveh ) );
    nand3_1 \I1/high/U1669/Und  ( .x(\I1/high/U1669/nd ), .a(
        \I1/high/ctrlack_internal ), .b(\I1/high/drivel ), .c(\I1/high/driveh 
        ) );
    oa21_1 \I1/high/U1669/U1  ( .x(\I1/high/U1669/n2 ), .a(\I1/high/U1669/n2 ), 
        .b(\I1/high/U1669/nr ), .c(\I1/high/U1669/nd ) );
    inv_2 \I1/high/U1669/U3  ( .x(\I1/net20 ), .a(\I1/high/U1669/n2 ) );
    buf_2 U1 ( .x(n1), .a(\I0/net20 ) );
    buf_1 U2 ( .x(n2), .a(\I0/low/latch ) );
    buf_2 U3 ( .x(n3), .a(net17) );
    buf_1 U4 ( .x(n4), .a(\I0/high/latch ) );
    buf_2 U5 ( .x(n5), .a(\I1/net20 ) );
    buf_1 U6 ( .x(n6), .a(\I1/low/latch ) );
    buf_2 U7 ( .x(n7), .a(ctrlreq) );
    buf_1 U8 ( .x(n8), .a(\I1/high/latch ) );
endmodule


module chain_irdemux_32new_3 ( ctrlack, oh, ol, pullreq, pull_h, pull_l, 
    pullcd, reset, ctrlreq );
output [31:0] oh;
output [31:0] ol;
input  [7:0] pull_h;
input  [7:0] pull_l;
input  pullcd, reset, ctrlreq;
output ctrlack, pullreq;
    wire net30, net31, net17, \I0/net20 , \I0/net33 , \I0/net32 , 
        \I0/low/drivel , \I0/low/driveh , \I0/low/localcd , \I0/low/ncd[7] , 
        \I0/low/ncd[6] , \I0/low/ncd[5] , \I0/low/ncd[4] , \I0/low/ncd[3] , 
        \I0/low/ncd[2] , \I0/low/ncd[1] , \I0/low/ncd[0] , \I0/low/ba , 
        \I0/low/latch , \I0/low/acb , \I0/low/ctrlack_internal , 
        \I0/low/nlocalcd , \I0/low/U4/U28/U1/clr , \I0/low/U4/U28/U1/set , 
        \I0/low/U1/Z , \I0/low/U1664/y[0] , \I0/low/U1664/y[1] , 
        \I0/low/U1664/x[1] , \I0/low/U1664/x[3] , \I0/low/U1664/x[2] , 
        \I0/low/U1664/x[0] , \I0/low/U1664/U28/Z , \I0/low/U1664/U32/Z , 
        \I0/low/U1664/U29/Z , \I0/low/U1664/U33/Z , \I0/low/U1664/U30/Z , 
        \I0/low/U1664/U31/Z , \I0/low/U1664/U37/Z , \I0/low/U1669/nr , 
        \I0/low/U1669/nd , \I0/low/U1669/n2 , \I0/high/drivel , 
        \I0/high/driveh , \I0/high/localcd , \I0/high/ncd[7] , 
        \I0/high/ncd[6] , \I0/high/ncd[5] , \I0/high/ncd[4] , \I0/high/ncd[3] , 
        \I0/high/ncd[2] , \I0/high/ncd[1] , \I0/high/ncd[0] , \I0/high/ba , 
        \I0/high/latch , \I0/high/acb , \I0/high/ctrlack_internal , 
        \I0/high/nlocalcd , \I0/high/U4/U28/U1/clr , \I0/high/U4/U28/U1/set , 
        \I0/high/U1/Z , \I0/high/U1664/y[0] , \I0/high/U1664/y[1] , 
        \I0/high/U1664/x[1] , \I0/high/U1664/x[3] , \I0/high/U1664/x[2] , 
        \I0/high/U1664/x[0] , \I0/high/U1664/U28/Z , \I0/high/U1664/U32/Z , 
        \I0/high/U1664/U29/Z , \I0/high/U1664/U33/Z , \I0/high/U1664/U30/Z , 
        \I0/high/U1664/U31/Z , \I0/high/U1664/U37/Z , \I0/high/U1669/nr , 
        \I0/high/U1669/nd , \I0/high/U1669/n2 , \I1/net20 , \I1/net33 , 
        \I1/net32 , \I1/low/drivel , \I1/low/driveh , \I1/low/localcd , 
        \I1/low/ncd[7] , \I1/low/ncd[6] , \I1/low/ncd[5] , \I1/low/ncd[4] , 
        \I1/low/ncd[3] , \I1/low/ncd[2] , \I1/low/ncd[1] , \I1/low/ncd[0] , 
        \I1/low/ba , \I1/low/latch , \I1/low/acb , \I1/low/ctrlack_internal , 
        \I1/low/nlocalcd , \I1/low/U4/U28/U1/clr , \I1/low/U4/U28/U1/set , 
        \I1/low/U1/Z , \I1/low/U1664/y[0] , \I1/low/U1664/y[1] , 
        \I1/low/U1664/x[1] , \I1/low/U1664/x[3] , \I1/low/U1664/x[2] , 
        \I1/low/U1664/x[0] , \I1/low/U1664/U28/Z , \I1/low/U1664/U32/Z , 
        \I1/low/U1664/U29/Z , \I1/low/U1664/U33/Z , \I1/low/U1664/U30/Z , 
        \I1/low/U1664/U31/Z , \I1/low/U1664/U37/Z , \I1/low/U1669/nr , 
        \I1/low/U1669/nd , \I1/low/U1669/n2 , \I1/high/localcd , 
        \I1/high/ncd[7] , \I1/high/ncd[6] , \I1/high/ncd[5] , \I1/high/ncd[4] , 
        \I1/high/ncd[3] , \I1/high/ncd[2] , \I1/high/ncd[1] , \I1/high/ncd[0] , 
        \I1/high/ba , \I1/high/latch , \I1/high/acb , 
        \I1/high/ctrlack_internal , \I1/high/nlocalcd , 
        \I1/high/U4/U28/U1/clr , \I1/high/U4/U28/U1/set , \I1/high/U1/Z , 
        \I1/high/U1664/y[0] , \I1/high/U1664/y[1] , \I1/high/U1664/x[1] , 
        \I1/high/U1664/x[3] , \I1/high/U1664/x[2] , \I1/high/U1664/x[0] , 
        \I1/high/U1664/U28/Z , \I1/high/U1664/U32/Z , \I1/high/U1664/U29/Z , 
        \I1/high/U1664/U33/Z , \I1/high/U1664/U30/Z , \I1/high/U1664/U31/Z , 
        \I1/high/U1664/U37/Z , \I1/high/U1669/nr , \I1/high/U1669/nd , 
        \I1/high/U1669/n2 , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
    nand2_1 \U3/U5  ( .x(pullreq), .a(net30), .b(net31) );
    nor2_1 \I0/U3/U5  ( .x(net30), .a(\I0/net32 ), .b(\I0/net33 ) );
    buf_2 \I0/low/U1653  ( .x(\I0/low/latch ), .a(\I0/net32 ) );
    nor2_1 \I0/low/U264/U5  ( .x(\I0/low/nlocalcd ), .a(reset), .b(
        \I0/low/localcd ) );
    nor2_1 \I0/low/U1659_0_/U5  ( .x(\I0/low/ncd[0] ), .a(ol[0]), .b(oh[0]) );
    nor2_1 \I0/low/U1659_1_/U5  ( .x(\I0/low/ncd[1] ), .a(ol[1]), .b(oh[1]) );
    nor2_1 \I0/low/U1659_2_/U5  ( .x(\I0/low/ncd[2] ), .a(ol[2]), .b(oh[2]) );
    nor2_1 \I0/low/U1659_3_/U5  ( .x(\I0/low/ncd[3] ), .a(ol[3]), .b(oh[3]) );
    nor2_1 \I0/low/U1659_4_/U5  ( .x(\I0/low/ncd[4] ), .a(ol[4]), .b(oh[4]) );
    nor2_1 \I0/low/U1659_5_/U5  ( .x(\I0/low/ncd[5] ), .a(ol[5]), .b(oh[5]) );
    nor2_1 \I0/low/U1659_6_/U5  ( .x(\I0/low/ncd[6] ), .a(ol[6]), .b(oh[6]) );
    nor2_1 \I0/low/U1659_7_/U5  ( .x(\I0/low/ncd[7] ), .a(ol[7]), .b(oh[7]) );
    nor2_1 \I0/low/U3/U5  ( .x(\I0/low/ctrlack_internal ), .a(\I0/low/acb ), 
        .b(\I0/low/ba ) );
    buf_2 \I0/low/U1665/U7  ( .x(\I0/low/driveh ), .a(\I0/net20 ) );
    buf_2 \I0/low/U1666/U7  ( .x(\I0/low/drivel ), .a(\I0/net20 ) );
    ao23_1 \I0/low/U1658_0_/U21/U1/U1  ( .x(ol[0]), .a(\I0/low/driveh ), .b(ol
        [0]), .c(n1), .d(pull_l[0]), .e(n2) );
    ao23_1 \I0/low/U1658_1_/U21/U1/U1  ( .x(ol[1]), .a(\I0/low/drivel ), .b(ol
        [1]), .c(\I0/low/driveh ), .d(pull_l[1]), .e(n2) );
    ao23_1 \I0/low/U1658_2_/U21/U1/U1  ( .x(ol[2]), .a(\I0/low/drivel ), .b(ol
        [2]), .c(\I0/low/driveh ), .d(pull_l[2]), .e(n2) );
    ao23_1 \I0/low/U1658_3_/U21/U1/U1  ( .x(ol[3]), .a(\I0/low/driveh ), .b(ol
        [3]), .c(\I0/low/drivel ), .d(pull_l[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_4_/U21/U1/U1  ( .x(ol[4]), .a(n1), .b(ol[4]), .c(
        \I0/low/drivel ), .d(pull_l[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_5_/U21/U1/U1  ( .x(ol[5]), .a(\I0/low/driveh ), .b(ol
        [5]), .c(n1), .d(pull_l[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_6_/U21/U1/U1  ( .x(ol[6]), .a(\I0/low/drivel ), .b(ol
        [6]), .c(\I0/low/driveh ), .d(pull_l[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_7_/U21/U1/U1  ( .x(ol[7]), .a(n1), .b(ol[7]), .c(n1), 
        .d(pull_l[7]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_0_/U21/U1/U1  ( .x(oh[0]), .a(\I0/low/driveh ), .b(oh
        [0]), .c(n1), .d(pull_h[0]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_1_/U21/U1/U1  ( .x(oh[1]), .a(n1), .b(oh[1]), .c(
        \I0/low/drivel ), .d(pull_h[1]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_2_/U21/U1/U1  ( .x(oh[2]), .a(\I0/low/drivel ), .b(oh
        [2]), .c(\I0/low/drivel ), .d(pull_h[2]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_3_/U21/U1/U1  ( .x(oh[3]), .a(n1), .b(oh[3]), .c(
        \I0/low/driveh ), .d(pull_h[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_4_/U21/U1/U1  ( .x(oh[4]), .a(n1), .b(oh[4]), .c(n1), 
        .d(pull_h[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_5_/U21/U1/U1  ( .x(oh[5]), .a(\I0/low/drivel ), .b(oh
        [5]), .c(n1), .d(pull_h[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_6_/U21/U1/U1  ( .x(oh[6]), .a(\I0/low/drivel ), .b(oh
        [6]), .c(\I0/low/driveh ), .d(pull_h[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_7_/U21/U1/U1  ( .x(oh[7]), .a(\I0/low/driveh ), .b(oh
        [7]), .c(\I0/low/drivel ), .d(pull_h[7]), .e(\I0/low/latch ) );
    aoai211_1 \I0/low/U4/U28/U1/U1  ( .x(\I0/low/U4/U28/U1/clr ), .a(
        \I0/net20 ), .b(\I0/low/acb ), .c(\I0/low/nlocalcd ), .d(\I0/net32 )
         );
    nand3_1 \I0/low/U4/U28/U1/U2  ( .x(\I0/low/U4/U28/U1/set ), .a(
        \I0/low/nlocalcd ), .b(\I0/net20 ), .c(\I0/low/acb ) );
    nand2_2 \I0/low/U4/U28/U1/U3  ( .x(\I0/net32 ), .a(\I0/low/U4/U28/U1/clr ), 
        .b(\I0/low/U4/U28/U1/set ) );
    oai21_1 \I0/low/U1/U30/U1/U1  ( .x(\I0/low/acb ), .a(\I0/low/U1/Z ), .b(
        \I0/low/ba ), .c(\I0/net20 ) );
    inv_1 \I0/low/U1/U30/U1/U2  ( .x(\I0/low/U1/Z ), .a(\I0/low/acb ) );
    ao222_1 \I0/low/U5/U18/U1/U1  ( .x(\I0/low/ba ), .a(\I0/low/latch ), .b(
        pullcd), .c(\I0/low/latch ), .d(\I0/low/ba ), .e(pullcd), .f(
        \I0/low/ba ) );
    aoi222_1 \I0/low/U1664/U28/U30/U1  ( .x(\I0/low/U1664/x[3] ), .a(
        \I0/low/ncd[7] ), .b(\I0/low/ncd[6] ), .c(\I0/low/ncd[7] ), .d(
        \I0/low/U1664/U28/Z ), .e(\I0/low/ncd[6] ), .f(\I0/low/U1664/U28/Z )
         );
    inv_1 \I0/low/U1664/U28/U30/Uinv  ( .x(\I0/low/U1664/U28/Z ), .a(
        \I0/low/U1664/x[3] ) );
    aoi222_1 \I0/low/U1664/U32/U30/U1  ( .x(\I0/low/U1664/x[0] ), .a(
        \I0/low/ncd[1] ), .b(\I0/low/ncd[0] ), .c(\I0/low/ncd[1] ), .d(
        \I0/low/U1664/U32/Z ), .e(\I0/low/ncd[0] ), .f(\I0/low/U1664/U32/Z )
         );
    inv_1 \I0/low/U1664/U32/U30/Uinv  ( .x(\I0/low/U1664/U32/Z ), .a(
        \I0/low/U1664/x[0] ) );
    aoi222_1 \I0/low/U1664/U29/U30/U1  ( .x(\I0/low/U1664/x[2] ), .a(
        \I0/low/ncd[5] ), .b(\I0/low/ncd[4] ), .c(\I0/low/ncd[5] ), .d(
        \I0/low/U1664/U29/Z ), .e(\I0/low/ncd[4] ), .f(\I0/low/U1664/U29/Z )
         );
    inv_1 \I0/low/U1664/U29/U30/Uinv  ( .x(\I0/low/U1664/U29/Z ), .a(
        \I0/low/U1664/x[2] ) );
    aoi222_1 \I0/low/U1664/U33/U30/U1  ( .x(\I0/low/U1664/y[0] ), .a(
        \I0/low/U1664/x[1] ), .b(\I0/low/U1664/x[0] ), .c(\I0/low/U1664/x[1] ), 
        .d(\I0/low/U1664/U33/Z ), .e(\I0/low/U1664/x[0] ), .f(
        \I0/low/U1664/U33/Z ) );
    inv_1 \I0/low/U1664/U33/U30/Uinv  ( .x(\I0/low/U1664/U33/Z ), .a(
        \I0/low/U1664/y[0] ) );
    aoi222_1 \I0/low/U1664/U30/U30/U1  ( .x(\I0/low/U1664/y[1] ), .a(
        \I0/low/U1664/x[3] ), .b(\I0/low/U1664/x[2] ), .c(\I0/low/U1664/x[3] ), 
        .d(\I0/low/U1664/U30/Z ), .e(\I0/low/U1664/x[2] ), .f(
        \I0/low/U1664/U30/Z ) );
    inv_1 \I0/low/U1664/U30/U30/Uinv  ( .x(\I0/low/U1664/U30/Z ), .a(
        \I0/low/U1664/y[1] ) );
    aoi222_1 \I0/low/U1664/U31/U30/U1  ( .x(\I0/low/U1664/x[1] ), .a(
        \I0/low/ncd[3] ), .b(\I0/low/ncd[2] ), .c(\I0/low/ncd[3] ), .d(
        \I0/low/U1664/U31/Z ), .e(\I0/low/ncd[2] ), .f(\I0/low/U1664/U31/Z )
         );
    inv_1 \I0/low/U1664/U31/U30/Uinv  ( .x(\I0/low/U1664/U31/Z ), .a(
        \I0/low/U1664/x[1] ) );
    aoi222_1 \I0/low/U1664/U37/U30/U1  ( .x(\I0/low/localcd ), .a(
        \I0/low/U1664/y[0] ), .b(\I0/low/U1664/y[1] ), .c(\I0/low/U1664/y[0] ), 
        .d(\I0/low/U1664/U37/Z ), .e(\I0/low/U1664/y[1] ), .f(
        \I0/low/U1664/U37/Z ) );
    inv_1 \I0/low/U1664/U37/U30/Uinv  ( .x(\I0/low/U1664/U37/Z ), .a(
        \I0/low/localcd ) );
    nor3_1 \I0/low/U1669/Unr  ( .x(\I0/low/U1669/nr ), .a(
        \I0/low/ctrlack_internal ), .b(n1), .c(\I0/low/driveh ) );
    nand3_1 \I0/low/U1669/Und  ( .x(\I0/low/U1669/nd ), .a(
        \I0/low/ctrlack_internal ), .b(\I0/low/drivel ), .c(\I0/low/driveh )
         );
    oa21_1 \I0/low/U1669/U1  ( .x(\I0/low/U1669/n2 ), .a(\I0/low/U1669/n2 ), 
        .b(\I0/low/U1669/nr ), .c(\I0/low/U1669/nd ) );
    inv_2 \I0/low/U1669/U3  ( .x(ctrlack), .a(\I0/low/U1669/n2 ) );
    buf_2 \I0/high/U1653  ( .x(\I0/high/latch ), .a(\I0/net33 ) );
    nor2_1 \I0/high/U264/U5  ( .x(\I0/high/nlocalcd ), .a(reset), .b(
        \I0/high/localcd ) );
    nor2_1 \I0/high/U1659_0_/U5  ( .x(\I0/high/ncd[0] ), .a(ol[8]), .b(oh[8])
         );
    nor2_1 \I0/high/U1659_1_/U5  ( .x(\I0/high/ncd[1] ), .a(ol[9]), .b(oh[9])
         );
    nor2_1 \I0/high/U1659_2_/U5  ( .x(\I0/high/ncd[2] ), .a(ol[10]), .b(oh[10]
        ) );
    nor2_1 \I0/high/U1659_3_/U5  ( .x(\I0/high/ncd[3] ), .a(ol[11]), .b(oh[11]
        ) );
    nor2_1 \I0/high/U1659_4_/U5  ( .x(\I0/high/ncd[4] ), .a(ol[12]), .b(oh[12]
        ) );
    nor2_1 \I0/high/U1659_5_/U5  ( .x(\I0/high/ncd[5] ), .a(ol[13]), .b(oh[13]
        ) );
    nor2_1 \I0/high/U1659_6_/U5  ( .x(\I0/high/ncd[6] ), .a(ol[14]), .b(oh[14]
        ) );
    nor2_1 \I0/high/U1659_7_/U5  ( .x(\I0/high/ncd[7] ), .a(ol[15]), .b(oh[15]
        ) );
    nor2_1 \I0/high/U3/U5  ( .x(\I0/high/ctrlack_internal ), .a(\I0/high/acb ), 
        .b(\I0/high/ba ) );
    buf_2 \I0/high/U1665/U7  ( .x(\I0/high/driveh ), .a(net17) );
    buf_2 \I0/high/U1666/U7  ( .x(\I0/high/drivel ), .a(net17) );
    ao23_1 \I0/high/U1658_0_/U21/U1/U1  ( .x(ol[8]), .a(\I0/high/driveh ), .b(
        ol[8]), .c(n3), .d(pull_l[0]), .e(n4) );
    ao23_1 \I0/high/U1658_1_/U21/U1/U1  ( .x(ol[9]), .a(\I0/high/drivel ), .b(
        ol[9]), .c(\I0/high/driveh ), .d(pull_l[1]), .e(n4) );
    ao23_1 \I0/high/U1658_2_/U21/U1/U1  ( .x(ol[10]), .a(\I0/high/drivel ), 
        .b(ol[10]), .c(\I0/high/driveh ), .d(pull_l[2]), .e(n4) );
    ao23_1 \I0/high/U1658_3_/U21/U1/U1  ( .x(ol[11]), .a(\I0/high/driveh ), 
        .b(ol[11]), .c(\I0/high/drivel ), .d(pull_l[3]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_4_/U21/U1/U1  ( .x(ol[12]), .a(n3), .b(ol[12]), .c(
        \I0/high/drivel ), .d(pull_l[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_5_/U21/U1/U1  ( .x(ol[13]), .a(\I0/high/driveh ), 
        .b(ol[13]), .c(n3), .d(pull_l[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_6_/U21/U1/U1  ( .x(ol[14]), .a(\I0/high/drivel ), 
        .b(ol[14]), .c(\I0/high/driveh ), .d(pull_l[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_7_/U21/U1/U1  ( .x(ol[15]), .a(n3), .b(ol[15]), .c(
        n3), .d(pull_l[7]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_0_/U21/U1/U1  ( .x(oh[8]), .a(\I0/high/driveh ), .b(
        oh[8]), .c(n3), .d(pull_h[0]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_1_/U21/U1/U1  ( .x(oh[9]), .a(n3), .b(oh[9]), .c(
        \I0/high/drivel ), .d(pull_h[1]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_2_/U21/U1/U1  ( .x(oh[10]), .a(\I0/high/drivel ), 
        .b(oh[10]), .c(\I0/high/drivel ), .d(pull_h[2]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_3_/U21/U1/U1  ( .x(oh[11]), .a(n3), .b(oh[11]), .c(
        \I0/high/driveh ), .d(pull_h[3]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_4_/U21/U1/U1  ( .x(oh[12]), .a(n3), .b(oh[12]), .c(
        n3), .d(pull_h[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_5_/U21/U1/U1  ( .x(oh[13]), .a(\I0/high/drivel ), 
        .b(oh[13]), .c(n3), .d(pull_h[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_6_/U21/U1/U1  ( .x(oh[14]), .a(\I0/high/drivel ), 
        .b(oh[14]), .c(\I0/high/driveh ), .d(pull_h[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_7_/U21/U1/U1  ( .x(oh[15]), .a(\I0/high/driveh ), 
        .b(oh[15]), .c(\I0/high/drivel ), .d(pull_h[7]), .e(\I0/high/latch )
         );
    aoai211_1 \I0/high/U4/U28/U1/U1  ( .x(\I0/high/U4/U28/U1/clr ), .a(net17), 
        .b(\I0/high/acb ), .c(\I0/high/nlocalcd ), .d(\I0/net33 ) );
    nand3_1 \I0/high/U4/U28/U1/U2  ( .x(\I0/high/U4/U28/U1/set ), .a(
        \I0/high/nlocalcd ), .b(net17), .c(\I0/high/acb ) );
    nand2_2 \I0/high/U4/U28/U1/U3  ( .x(\I0/net33 ), .a(
        \I0/high/U4/U28/U1/clr ), .b(\I0/high/U4/U28/U1/set ) );
    oai21_1 \I0/high/U1/U30/U1/U1  ( .x(\I0/high/acb ), .a(\I0/high/U1/Z ), 
        .b(\I0/high/ba ), .c(net17) );
    inv_1 \I0/high/U1/U30/U1/U2  ( .x(\I0/high/U1/Z ), .a(\I0/high/acb ) );
    ao222_1 \I0/high/U5/U18/U1/U1  ( .x(\I0/high/ba ), .a(\I0/high/latch ), 
        .b(pullcd), .c(\I0/high/latch ), .d(\I0/high/ba ), .e(pullcd), .f(
        \I0/high/ba ) );
    aoi222_1 \I0/high/U1664/U28/U30/U1  ( .x(\I0/high/U1664/x[3] ), .a(
        \I0/high/ncd[7] ), .b(\I0/high/ncd[6] ), .c(\I0/high/ncd[7] ), .d(
        \I0/high/U1664/U28/Z ), .e(\I0/high/ncd[6] ), .f(\I0/high/U1664/U28/Z 
        ) );
    inv_1 \I0/high/U1664/U28/U30/Uinv  ( .x(\I0/high/U1664/U28/Z ), .a(
        \I0/high/U1664/x[3] ) );
    aoi222_1 \I0/high/U1664/U32/U30/U1  ( .x(\I0/high/U1664/x[0] ), .a(
        \I0/high/ncd[1] ), .b(\I0/high/ncd[0] ), .c(\I0/high/ncd[1] ), .d(
        \I0/high/U1664/U32/Z ), .e(\I0/high/ncd[0] ), .f(\I0/high/U1664/U32/Z 
        ) );
    inv_1 \I0/high/U1664/U32/U30/Uinv  ( .x(\I0/high/U1664/U32/Z ), .a(
        \I0/high/U1664/x[0] ) );
    aoi222_1 \I0/high/U1664/U29/U30/U1  ( .x(\I0/high/U1664/x[2] ), .a(
        \I0/high/ncd[5] ), .b(\I0/high/ncd[4] ), .c(\I0/high/ncd[5] ), .d(
        \I0/high/U1664/U29/Z ), .e(\I0/high/ncd[4] ), .f(\I0/high/U1664/U29/Z 
        ) );
    inv_1 \I0/high/U1664/U29/U30/Uinv  ( .x(\I0/high/U1664/U29/Z ), .a(
        \I0/high/U1664/x[2] ) );
    aoi222_1 \I0/high/U1664/U33/U30/U1  ( .x(\I0/high/U1664/y[0] ), .a(
        \I0/high/U1664/x[1] ), .b(\I0/high/U1664/x[0] ), .c(
        \I0/high/U1664/x[1] ), .d(\I0/high/U1664/U33/Z ), .e(
        \I0/high/U1664/x[0] ), .f(\I0/high/U1664/U33/Z ) );
    inv_1 \I0/high/U1664/U33/U30/Uinv  ( .x(\I0/high/U1664/U33/Z ), .a(
        \I0/high/U1664/y[0] ) );
    aoi222_1 \I0/high/U1664/U30/U30/U1  ( .x(\I0/high/U1664/y[1] ), .a(
        \I0/high/U1664/x[3] ), .b(\I0/high/U1664/x[2] ), .c(
        \I0/high/U1664/x[3] ), .d(\I0/high/U1664/U30/Z ), .e(
        \I0/high/U1664/x[2] ), .f(\I0/high/U1664/U30/Z ) );
    inv_1 \I0/high/U1664/U30/U30/Uinv  ( .x(\I0/high/U1664/U30/Z ), .a(
        \I0/high/U1664/y[1] ) );
    aoi222_1 \I0/high/U1664/U31/U30/U1  ( .x(\I0/high/U1664/x[1] ), .a(
        \I0/high/ncd[3] ), .b(\I0/high/ncd[2] ), .c(\I0/high/ncd[3] ), .d(
        \I0/high/U1664/U31/Z ), .e(\I0/high/ncd[2] ), .f(\I0/high/U1664/U31/Z 
        ) );
    inv_1 \I0/high/U1664/U31/U30/Uinv  ( .x(\I0/high/U1664/U31/Z ), .a(
        \I0/high/U1664/x[1] ) );
    aoi222_1 \I0/high/U1664/U37/U30/U1  ( .x(\I0/high/localcd ), .a(
        \I0/high/U1664/y[0] ), .b(\I0/high/U1664/y[1] ), .c(
        \I0/high/U1664/y[0] ), .d(\I0/high/U1664/U37/Z ), .e(
        \I0/high/U1664/y[1] ), .f(\I0/high/U1664/U37/Z ) );
    inv_1 \I0/high/U1664/U37/U30/Uinv  ( .x(\I0/high/U1664/U37/Z ), .a(
        \I0/high/localcd ) );
    nor3_1 \I0/high/U1669/Unr  ( .x(\I0/high/U1669/nr ), .a(
        \I0/high/ctrlack_internal ), .b(n3), .c(\I0/high/driveh ) );
    nand3_1 \I0/high/U1669/Und  ( .x(\I0/high/U1669/nd ), .a(
        \I0/high/ctrlack_internal ), .b(\I0/high/drivel ), .c(\I0/high/driveh 
        ) );
    oa21_1 \I0/high/U1669/U1  ( .x(\I0/high/U1669/n2 ), .a(\I0/high/U1669/n2 ), 
        .b(\I0/high/U1669/nr ), .c(\I0/high/U1669/nd ) );
    inv_2 \I0/high/U1669/U3  ( .x(\I0/net20 ), .a(\I0/high/U1669/n2 ) );
    nor2_1 \I1/U3/U5  ( .x(net31), .a(\I1/net32 ), .b(\I1/net33 ) );
    buf_2 \I1/low/U1653  ( .x(\I1/low/latch ), .a(\I1/net32 ) );
    nor2_1 \I1/low/U264/U5  ( .x(\I1/low/nlocalcd ), .a(reset), .b(
        \I1/low/localcd ) );
    nor2_1 \I1/low/U1659_0_/U5  ( .x(\I1/low/ncd[0] ), .a(ol[16]), .b(oh[16])
         );
    nor2_1 \I1/low/U1659_1_/U5  ( .x(\I1/low/ncd[1] ), .a(ol[17]), .b(oh[17])
         );
    nor2_1 \I1/low/U1659_2_/U5  ( .x(\I1/low/ncd[2] ), .a(ol[18]), .b(oh[18])
         );
    nor2_1 \I1/low/U1659_3_/U5  ( .x(\I1/low/ncd[3] ), .a(ol[19]), .b(oh[19])
         );
    nor2_1 \I1/low/U1659_4_/U5  ( .x(\I1/low/ncd[4] ), .a(ol[20]), .b(oh[20])
         );
    nor2_1 \I1/low/U1659_5_/U5  ( .x(\I1/low/ncd[5] ), .a(ol[21]), .b(oh[21])
         );
    nor2_1 \I1/low/U1659_6_/U5  ( .x(\I1/low/ncd[6] ), .a(ol[22]), .b(oh[22])
         );
    nor2_1 \I1/low/U1659_7_/U5  ( .x(\I1/low/ncd[7] ), .a(ol[23]), .b(oh[23])
         );
    nor2_1 \I1/low/U3/U5  ( .x(\I1/low/ctrlack_internal ), .a(\I1/low/acb ), 
        .b(\I1/low/ba ) );
    buf_2 \I1/low/U1665/U7  ( .x(\I1/low/driveh ), .a(\I1/net20 ) );
    buf_2 \I1/low/U1666/U7  ( .x(\I1/low/drivel ), .a(\I1/net20 ) );
    ao23_1 \I1/low/U1658_0_/U21/U1/U1  ( .x(ol[16]), .a(\I1/low/drivel ), .b(
        ol[16]), .c(n5), .d(pull_l[0]), .e(n6) );
    ao23_1 \I1/low/U1658_1_/U21/U1/U1  ( .x(ol[17]), .a(\I1/low/driveh ), .b(
        ol[17]), .c(n5), .d(pull_l[1]), .e(n6) );
    ao23_1 \I1/low/U1658_2_/U21/U1/U1  ( .x(ol[18]), .a(\I1/low/drivel ), .b(
        ol[18]), .c(\I1/low/driveh ), .d(pull_l[2]), .e(n6) );
    ao23_1 \I1/low/U1658_3_/U21/U1/U1  ( .x(ol[19]), .a(n5), .b(ol[19]), .c(
        \I1/low/driveh ), .d(pull_l[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_4_/U21/U1/U1  ( .x(ol[20]), .a(\I1/low/driveh ), .b(
        ol[20]), .c(\I1/low/drivel ), .d(pull_l[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_5_/U21/U1/U1  ( .x(ol[21]), .a(n5), .b(ol[21]), .c(
        \I1/low/drivel ), .d(pull_l[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_6_/U21/U1/U1  ( .x(ol[22]), .a(\I1/low/driveh ), .b(
        ol[22]), .c(n5), .d(pull_l[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_7_/U21/U1/U1  ( .x(ol[23]), .a(\I1/low/drivel ), .b(
        ol[23]), .c(\I1/low/driveh ), .d(pull_l[7]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_0_/U21/U1/U1  ( .x(oh[16]), .a(\I1/low/driveh ), .b(
        oh[16]), .c(\I1/low/drivel ), .d(pull_h[0]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_1_/U21/U1/U1  ( .x(oh[17]), .a(\I1/low/drivel ), .b(
        oh[17]), .c(n5), .d(pull_h[1]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_2_/U21/U1/U1  ( .x(oh[18]), .a(\I1/low/drivel ), .b(
        oh[18]), .c(\I1/low/driveh ), .d(pull_h[2]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_3_/U21/U1/U1  ( .x(oh[19]), .a(n5), .b(oh[19]), .c(n5
        ), .d(pull_h[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_4_/U21/U1/U1  ( .x(oh[20]), .a(n5), .b(oh[20]), .c(n5
        ), .d(pull_h[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_5_/U21/U1/U1  ( .x(oh[21]), .a(\I1/low/drivel ), .b(
        oh[21]), .c(\I1/low/driveh ), .d(pull_h[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_6_/U21/U1/U1  ( .x(oh[22]), .a(n5), .b(oh[22]), .c(
        \I1/low/drivel ), .d(pull_h[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_7_/U21/U1/U1  ( .x(oh[23]), .a(\I1/low/driveh ), .b(
        oh[23]), .c(\I1/low/drivel ), .d(pull_h[7]), .e(\I1/low/latch ) );
    aoai211_1 \I1/low/U4/U28/U1/U1  ( .x(\I1/low/U4/U28/U1/clr ), .a(
        \I1/net20 ), .b(\I1/low/acb ), .c(\I1/low/nlocalcd ), .d(\I1/net32 )
         );
    nand3_1 \I1/low/U4/U28/U1/U2  ( .x(\I1/low/U4/U28/U1/set ), .a(
        \I1/low/nlocalcd ), .b(\I1/net20 ), .c(\I1/low/acb ) );
    nand2_2 \I1/low/U4/U28/U1/U3  ( .x(\I1/net32 ), .a(\I1/low/U4/U28/U1/clr ), 
        .b(\I1/low/U4/U28/U1/set ) );
    oai21_1 \I1/low/U1/U30/U1/U1  ( .x(\I1/low/acb ), .a(\I1/low/U1/Z ), .b(
        \I1/low/ba ), .c(\I1/net20 ) );
    inv_1 \I1/low/U1/U30/U1/U2  ( .x(\I1/low/U1/Z ), .a(\I1/low/acb ) );
    ao222_1 \I1/low/U5/U18/U1/U1  ( .x(\I1/low/ba ), .a(\I1/low/latch ), .b(
        pullcd), .c(\I1/low/latch ), .d(\I1/low/ba ), .e(pullcd), .f(
        \I1/low/ba ) );
    aoi222_1 \I1/low/U1664/U28/U30/U1  ( .x(\I1/low/U1664/x[3] ), .a(
        \I1/low/ncd[7] ), .b(\I1/low/ncd[6] ), .c(\I1/low/ncd[7] ), .d(
        \I1/low/U1664/U28/Z ), .e(\I1/low/ncd[6] ), .f(\I1/low/U1664/U28/Z )
         );
    inv_1 \I1/low/U1664/U28/U30/Uinv  ( .x(\I1/low/U1664/U28/Z ), .a(
        \I1/low/U1664/x[3] ) );
    aoi222_1 \I1/low/U1664/U32/U30/U1  ( .x(\I1/low/U1664/x[0] ), .a(
        \I1/low/ncd[1] ), .b(\I1/low/ncd[0] ), .c(\I1/low/ncd[1] ), .d(
        \I1/low/U1664/U32/Z ), .e(\I1/low/ncd[0] ), .f(\I1/low/U1664/U32/Z )
         );
    inv_1 \I1/low/U1664/U32/U30/Uinv  ( .x(\I1/low/U1664/U32/Z ), .a(
        \I1/low/U1664/x[0] ) );
    aoi222_1 \I1/low/U1664/U29/U30/U1  ( .x(\I1/low/U1664/x[2] ), .a(
        \I1/low/ncd[5] ), .b(\I1/low/ncd[4] ), .c(\I1/low/ncd[5] ), .d(
        \I1/low/U1664/U29/Z ), .e(\I1/low/ncd[4] ), .f(\I1/low/U1664/U29/Z )
         );
    inv_1 \I1/low/U1664/U29/U30/Uinv  ( .x(\I1/low/U1664/U29/Z ), .a(
        \I1/low/U1664/x[2] ) );
    aoi222_1 \I1/low/U1664/U33/U30/U1  ( .x(\I1/low/U1664/y[0] ), .a(
        \I1/low/U1664/x[1] ), .b(\I1/low/U1664/x[0] ), .c(\I1/low/U1664/x[1] ), 
        .d(\I1/low/U1664/U33/Z ), .e(\I1/low/U1664/x[0] ), .f(
        \I1/low/U1664/U33/Z ) );
    inv_1 \I1/low/U1664/U33/U30/Uinv  ( .x(\I1/low/U1664/U33/Z ), .a(
        \I1/low/U1664/y[0] ) );
    aoi222_1 \I1/low/U1664/U30/U30/U1  ( .x(\I1/low/U1664/y[1] ), .a(
        \I1/low/U1664/x[3] ), .b(\I1/low/U1664/x[2] ), .c(\I1/low/U1664/x[3] ), 
        .d(\I1/low/U1664/U30/Z ), .e(\I1/low/U1664/x[2] ), .f(
        \I1/low/U1664/U30/Z ) );
    inv_1 \I1/low/U1664/U30/U30/Uinv  ( .x(\I1/low/U1664/U30/Z ), .a(
        \I1/low/U1664/y[1] ) );
    aoi222_1 \I1/low/U1664/U31/U30/U1  ( .x(\I1/low/U1664/x[1] ), .a(
        \I1/low/ncd[3] ), .b(\I1/low/ncd[2] ), .c(\I1/low/ncd[3] ), .d(
        \I1/low/U1664/U31/Z ), .e(\I1/low/ncd[2] ), .f(\I1/low/U1664/U31/Z )
         );
    inv_1 \I1/low/U1664/U31/U30/Uinv  ( .x(\I1/low/U1664/U31/Z ), .a(
        \I1/low/U1664/x[1] ) );
    aoi222_1 \I1/low/U1664/U37/U30/U1  ( .x(\I1/low/localcd ), .a(
        \I1/low/U1664/y[0] ), .b(\I1/low/U1664/y[1] ), .c(\I1/low/U1664/y[0] ), 
        .d(\I1/low/U1664/U37/Z ), .e(\I1/low/U1664/y[1] ), .f(
        \I1/low/U1664/U37/Z ) );
    inv_1 \I1/low/U1664/U37/U30/Uinv  ( .x(\I1/low/U1664/U37/Z ), .a(
        \I1/low/localcd ) );
    nor3_1 \I1/low/U1669/Unr  ( .x(\I1/low/U1669/nr ), .a(
        \I1/low/ctrlack_internal ), .b(n5), .c(\I1/low/driveh ) );
    nand3_1 \I1/low/U1669/Und  ( .x(\I1/low/U1669/nd ), .a(
        \I1/low/ctrlack_internal ), .b(\I1/low/drivel ), .c(\I1/low/driveh )
         );
    oa21_1 \I1/low/U1669/U1  ( .x(\I1/low/U1669/n2 ), .a(\I1/low/U1669/n2 ), 
        .b(\I1/low/U1669/nr ), .c(\I1/low/U1669/nd ) );
    inv_2 \I1/low/U1669/U3  ( .x(net17), .a(\I1/low/U1669/n2 ) );
    buf_2 \I1/high/U1653  ( .x(\I1/high/latch ), .a(\I1/net33 ) );
    nor2_1 \I1/high/U264/U5  ( .x(\I1/high/nlocalcd ), .a(reset), .b(
        \I1/high/localcd ) );
    nor2_1 \I1/high/U1659_0_/U5  ( .x(\I1/high/ncd[0] ), .a(ol[24]), .b(oh[24]
        ) );
    nor2_1 \I1/high/U1659_1_/U5  ( .x(\I1/high/ncd[1] ), .a(ol[25]), .b(oh[25]
        ) );
    nor2_1 \I1/high/U1659_2_/U5  ( .x(\I1/high/ncd[2] ), .a(ol[26]), .b(oh[26]
        ) );
    nor2_1 \I1/high/U1659_3_/U5  ( .x(\I1/high/ncd[3] ), .a(ol[27]), .b(oh[27]
        ) );
    nor2_1 \I1/high/U1659_4_/U5  ( .x(\I1/high/ncd[4] ), .a(ol[28]), .b(oh[28]
        ) );
    nor2_1 \I1/high/U1659_5_/U5  ( .x(\I1/high/ncd[5] ), .a(ol[29]), .b(oh[29]
        ) );
    nor2_1 \I1/high/U1659_6_/U5  ( .x(\I1/high/ncd[6] ), .a(ol[30]), .b(oh[30]
        ) );
    nor2_1 \I1/high/U1659_7_/U5  ( .x(\I1/high/ncd[7] ), .a(ol[31]), .b(oh[31]
        ) );
    nor2_1 \I1/high/U3/U5  ( .x(\I1/high/ctrlack_internal ), .a(\I1/high/acb ), 
        .b(\I1/high/ba ) );
    ao23_1 \I1/high/U1658_0_/U21/U1/U1  ( .x(ol[24]), .a(n7), .b(ol[24]), .c(
        n8), .d(pull_l[0]), .e(n12) );
    ao23_1 \I1/high/U1658_1_/U21/U1/U1  ( .x(ol[25]), .a(n7), .b(ol[25]), .c(
        n8), .d(pull_l[1]), .e(n12) );
    ao23_1 \I1/high/U1658_2_/U21/U1/U1  ( .x(ol[26]), .a(n7), .b(ol[26]), .c(
        n7), .d(pull_l[2]), .e(n12) );
    ao23_1 \I1/high/U1658_3_/U21/U1/U1  ( .x(ol[27]), .a(n7), .b(ol[27]), .c(
        n7), .d(pull_l[3]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_4_/U21/U1/U1  ( .x(ol[28]), .a(n7), .b(ol[28]), .c(
        n7), .d(pull_l[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_5_/U21/U1/U1  ( .x(ol[29]), .a(n7), .b(ol[29]), .c(
        n8), .d(pull_l[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_6_/U21/U1/U1  ( .x(ol[30]), .a(n7), .b(ol[30]), .c(
        n8), .d(pull_l[6]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_7_/U21/U1/U1  ( .x(ol[31]), .a(n7), .b(ol[31]), .c(
        n8), .d(pull_l[7]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_0_/U21/U1/U1  ( .x(oh[24]), .a(n10), .b(oh[24]), .c(
        n10), .d(pull_h[0]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_1_/U21/U1/U1  ( .x(oh[25]), .a(n10), .b(oh[25]), .c(
        n11), .d(pull_h[1]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_2_/U21/U1/U1  ( .x(oh[26]), .a(n10), .b(oh[26]), .c(
        n11), .d(pull_h[2]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_3_/U21/U1/U1  ( .x(oh[27]), .a(n10), .b(oh[27]), .c(
        n10), .d(pull_h[3]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_4_/U21/U1/U1  ( .x(oh[28]), .a(n10), .b(oh[28]), .c(
        n11), .d(pull_h[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_5_/U21/U1/U1  ( .x(oh[29]), .a(n10), .b(oh[29]), .c(
        n11), .d(pull_h[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_6_/U21/U1/U1  ( .x(oh[30]), .a(n10), .b(oh[30]), .c(
        n11), .d(pull_h[6]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_7_/U21/U1/U1  ( .x(oh[31]), .a(n10), .b(oh[31]), .c(
        n10), .d(pull_h[7]), .e(\I1/high/latch ) );
    aoai211_1 \I1/high/U4/U28/U1/U1  ( .x(\I1/high/U4/U28/U1/clr ), .a(ctrlreq
        ), .b(\I1/high/acb ), .c(\I1/high/nlocalcd ), .d(\I1/net33 ) );
    nand3_1 \I1/high/U4/U28/U1/U2  ( .x(\I1/high/U4/U28/U1/set ), .a(
        \I1/high/nlocalcd ), .b(ctrlreq), .c(\I1/high/acb ) );
    nand2_2 \I1/high/U4/U28/U1/U3  ( .x(\I1/net33 ), .a(
        \I1/high/U4/U28/U1/clr ), .b(\I1/high/U4/U28/U1/set ) );
    oai21_1 \I1/high/U1/U30/U1/U1  ( .x(\I1/high/acb ), .a(\I1/high/U1/Z ), 
        .b(\I1/high/ba ), .c(ctrlreq) );
    inv_1 \I1/high/U1/U30/U1/U2  ( .x(\I1/high/U1/Z ), .a(\I1/high/acb ) );
    ao222_1 \I1/high/U5/U18/U1/U1  ( .x(\I1/high/ba ), .a(\I1/high/latch ), 
        .b(pullcd), .c(\I1/high/latch ), .d(\I1/high/ba ), .e(pullcd), .f(
        \I1/high/ba ) );
    aoi222_1 \I1/high/U1664/U28/U30/U1  ( .x(\I1/high/U1664/x[3] ), .a(
        \I1/high/ncd[7] ), .b(\I1/high/ncd[6] ), .c(\I1/high/ncd[7] ), .d(
        \I1/high/U1664/U28/Z ), .e(\I1/high/ncd[6] ), .f(\I1/high/U1664/U28/Z 
        ) );
    inv_1 \I1/high/U1664/U28/U30/Uinv  ( .x(\I1/high/U1664/U28/Z ), .a(
        \I1/high/U1664/x[3] ) );
    aoi222_1 \I1/high/U1664/U32/U30/U1  ( .x(\I1/high/U1664/x[0] ), .a(
        \I1/high/ncd[1] ), .b(\I1/high/ncd[0] ), .c(\I1/high/ncd[1] ), .d(
        \I1/high/U1664/U32/Z ), .e(\I1/high/ncd[0] ), .f(\I1/high/U1664/U32/Z 
        ) );
    inv_1 \I1/high/U1664/U32/U30/Uinv  ( .x(\I1/high/U1664/U32/Z ), .a(
        \I1/high/U1664/x[0] ) );
    aoi222_1 \I1/high/U1664/U29/U30/U1  ( .x(\I1/high/U1664/x[2] ), .a(
        \I1/high/ncd[5] ), .b(\I1/high/ncd[4] ), .c(\I1/high/ncd[5] ), .d(
        \I1/high/U1664/U29/Z ), .e(\I1/high/ncd[4] ), .f(\I1/high/U1664/U29/Z 
        ) );
    inv_1 \I1/high/U1664/U29/U30/Uinv  ( .x(\I1/high/U1664/U29/Z ), .a(
        \I1/high/U1664/x[2] ) );
    aoi222_1 \I1/high/U1664/U33/U30/U1  ( .x(\I1/high/U1664/y[0] ), .a(
        \I1/high/U1664/x[1] ), .b(\I1/high/U1664/x[0] ), .c(
        \I1/high/U1664/x[1] ), .d(\I1/high/U1664/U33/Z ), .e(
        \I1/high/U1664/x[0] ), .f(\I1/high/U1664/U33/Z ) );
    inv_1 \I1/high/U1664/U33/U30/Uinv  ( .x(\I1/high/U1664/U33/Z ), .a(
        \I1/high/U1664/y[0] ) );
    aoi222_1 \I1/high/U1664/U30/U30/U1  ( .x(\I1/high/U1664/y[1] ), .a(
        \I1/high/U1664/x[3] ), .b(\I1/high/U1664/x[2] ), .c(
        \I1/high/U1664/x[3] ), .d(\I1/high/U1664/U30/Z ), .e(
        \I1/high/U1664/x[2] ), .f(\I1/high/U1664/U30/Z ) );
    inv_1 \I1/high/U1664/U30/U30/Uinv  ( .x(\I1/high/U1664/U30/Z ), .a(
        \I1/high/U1664/y[1] ) );
    aoi222_1 \I1/high/U1664/U31/U30/U1  ( .x(\I1/high/U1664/x[1] ), .a(
        \I1/high/ncd[3] ), .b(\I1/high/ncd[2] ), .c(\I1/high/ncd[3] ), .d(
        \I1/high/U1664/U31/Z ), .e(\I1/high/ncd[2] ), .f(\I1/high/U1664/U31/Z 
        ) );
    inv_1 \I1/high/U1664/U31/U30/Uinv  ( .x(\I1/high/U1664/U31/Z ), .a(
        \I1/high/U1664/x[1] ) );
    aoi222_1 \I1/high/U1664/U37/U30/U1  ( .x(\I1/high/localcd ), .a(
        \I1/high/U1664/y[0] ), .b(\I1/high/U1664/y[1] ), .c(
        \I1/high/U1664/y[0] ), .d(\I1/high/U1664/U37/Z ), .e(
        \I1/high/U1664/y[1] ), .f(\I1/high/U1664/U37/Z ) );
    inv_1 \I1/high/U1664/U37/U30/Uinv  ( .x(\I1/high/U1664/U37/Z ), .a(
        \I1/high/localcd ) );
    nor3_1 \I1/high/U1669/Unr  ( .x(\I1/high/U1669/nr ), .a(
        \I1/high/ctrlack_internal ), .b(n8), .c(n11) );
    nand3_1 \I1/high/U1669/Und  ( .x(\I1/high/U1669/nd ), .a(
        \I1/high/ctrlack_internal ), .b(n8), .c(n11) );
    oa21_1 \I1/high/U1669/U1  ( .x(\I1/high/U1669/n2 ), .a(\I1/high/U1669/n2 ), 
        .b(\I1/high/U1669/nr ), .c(\I1/high/U1669/nd ) );
    inv_2 \I1/high/U1669/U3  ( .x(\I1/net20 ), .a(\I1/high/U1669/n2 ) );
    buf_2 U1 ( .x(n1), .a(\I0/net20 ) );
    buf_1 U2 ( .x(n2), .a(\I0/low/latch ) );
    buf_2 U3 ( .x(n3), .a(net17) );
    buf_1 U4 ( .x(n4), .a(\I0/high/latch ) );
    buf_2 U5 ( .x(n5), .a(\I1/net20 ) );
    buf_1 U6 ( .x(n6), .a(\I1/low/latch ) );
    inv_2 U7 ( .x(n7), .a(n9) );
    inv_1 U8 ( .x(n8), .a(n9) );
    inv_0 U9 ( .x(n9), .a(ctrlreq) );
    inv_2 U10 ( .x(n10), .a(n9) );
    inv_1 U11 ( .x(n11), .a(n9) );
    buf_1 U12 ( .x(n12), .a(\I1/high/latch ) );
endmodule


module chain_fr2dr_byte_1 ( nia, oh, ol, i, nReset, noa );
output [7:0] oh;
output [7:0] ol;
input  [4:0] i;
input  nReset, noa;
output nia;
    wire eop, net135, nca, nbReset, ncla, \c[3] , \c[2] , \c[1] , \c[0] , 
        \cl[3] , \cl[2] , \cl[1] , \cl[0] , asel, bsel, asela, bsela, csel, 
        dsel, csela, dsela, esel, fsel, esela, fsela, naa, nda, \a[3] , \a[2] , 
        \a[1] , \a[0] , \d[3] , \d[2] , \d[1] , \d[0] , nba, nea, nfa, \b[3] , 
        \b[2] , \b[1] , \b[0] , \f[3] , \f[2] , \f[1] , \f[0] , \e[3] , \e[2] , 
        \e[1] , \e[0] , \U891/nack , \U891/acka , \U891/naack[0] , 
        \U891/naack[1] , \U891/iay , \U891/ackb , \U891/reset , \U891/neopack , 
        \U891/U1128/nb , \U891/U1128/na , \U891/U1118_0_/nr , 
        \U891/U1118_0_/nd , \U891/U1118_0_/n2 , \U891/U1118_1_/nr , 
        \U891/U1118_1_/nd , \U891/U1118_1_/n2 , \U891/U1118_2_/nr , 
        \U891/U1118_2_/nd , \U891/U1118_2_/n2 , \U891/U1118_3_/nr , 
        \U891/U1118_3_/nd , \U891/U1118_3_/n2 , \U891/U1117_0_/nr , 
        \U891/U1117_0_/nd , \U891/U1117_0_/n2 , \U891/U1117_1_/nr , 
        \U891/U1117_1_/nd , \U891/U1117_1_/n2 , \U891/U1117_2_/nr , 
        \U891/U1117_2_/nd , \U891/U1117_2_/n2 , \U891/U1117_3_/nr , 
        \U891/U1117_3_/nd , \U891/U1117_3_/n2 , \U886/nack , \U886/acka , 
        \U886/ackb , \U886/reset , \U886/U1128/nb , \U886/U1128/na , 
        \U886/U1127/n5 , \U886/U1127/n1 , \U886/U1127/n2 , \U886/U1127/n3 , 
        \U886/U1127/n4 , \U886/U1118_0_/nr , \U886/U1118_0_/nd , 
        \U886/U1118_0_/n2 , \U886/U1118_1_/nr , \U886/U1118_1_/nd , 
        \U886/U1118_1_/n2 , \U886/U1118_2_/nr , \U886/U1118_2_/nd , 
        \U886/U1118_2_/n2 , \U886/U1118_3_/nr , \U886/U1118_3_/nd , 
        \U886/U1118_3_/n2 , \U886/U1117_0_/nr , \U886/U1117_0_/nd , 
        \U886/U1117_0_/n2 , \U886/U1117_1_/nr , \U886/U1117_1_/nd , 
        \U886/U1117_1_/n2 , \U886/U1117_2_/nr , \U886/U1117_2_/nd , 
        \U886/U1117_2_/n2 , \U886/U1117_3_/nr , \U886/U1117_3_/nd , 
        \U886/U1117_3_/n2 , \U884/nack , \U884/acka , \U884/ackb , 
        \U884/reset , \U884/U1128/nb , \U884/U1128/na , \U884/U1127/n5 , 
        \U884/U1127/n1 , \U884/U1127/n2 , \U884/U1127/n3 , \U884/U1127/n4 , 
        \U884/U1118_0_/nr , \U884/U1118_0_/nd , \U884/U1118_0_/n2 , 
        \U884/U1118_1_/nr , \U884/U1118_1_/nd , \U884/U1118_1_/n2 , 
        \U884/U1118_2_/nr , \U884/U1118_2_/nd , \U884/U1118_2_/n2 , 
        \U884/U1118_3_/nr , \U884/U1118_3_/nd , \U884/U1118_3_/n2 , 
        \U884/U1117_0_/nr , \U884/U1117_0_/nd , \U884/U1117_0_/n2 , 
        \U884/U1117_1_/nr , \U884/U1117_1_/nd , \U884/U1117_1_/n2 , 
        \U884/U1117_2_/nr , \U884/U1117_2_/nd , \U884/U1117_2_/n2 , 
        \U884/U1117_3_/nr , \U884/U1117_3_/nd , \U884/U1117_3_/n2 , 
        \U888/naack , \U888/r , \U888/s , \U888/nback , \U888/reset , 
        \U887/naack , \U887/r , \U887/s , \U887/nback , \U887/reset , 
        \U885/naack , \U885/r , \U885/s , \U885/nback , \U885/reset , \U877/x , 
        \U877/y , \U877/reset , \U877/U590/U25/U1/clr , \U877/U590/U25/U1/ob , 
        \U877/U589/U25/U1/clr , \U877/U589/U25/U1/ob , \U877/U588/U25/U1/clr , 
        \U877/U588/U25/U1/ob , \U877/U591/U25/U1/clr , \U877/U591/U25/U1/ob , 
        \U876/x , \U876/y , \U876/reset , \U876/U590/U25/U1/clr , 
        \U876/U590/U25/U1/ob , \U876/U589/U25/U1/clr , \U876/U589/U25/U1/ob , 
        \U876/U588/U25/U1/clr , \U876/U588/U25/U1/ob , \U876/U591/U25/U1/clr , 
        \U876/U591/U25/U1/ob , \U2/x , \U2/y , \U2/reset , 
        \U2/U590/U25/U1/clr , \U2/U590/U25/U1/ob , \U2/U589/U25/U1/clr , 
        \U2/U589/U25/U1/ob , \U2/U588/U25/U1/clr , \U2/U588/U25/U1/ob , 
        \U2/U591/U25/U1/clr , \U2/U591/U25/U1/ob , \U1/x , \U1/y , \U1/reset , 
        \U1/U590/U25/U1/clr , \U1/U590/U25/U1/ob , \U1/U589/U25/U1/clr , 
        \U1/U589/U25/U1/ob , \U1/U588/U25/U1/clr , \U1/U588/U25/U1/ob , 
        \U1/U591/U25/U1/clr , \U1/U591/U25/U1/ob , \U881/nack[1] , 
        \U881/nack[0] , n1;
    buf_2 U897 ( .x(nbReset), .a(nReset) );
    and4_1 \U894/U12  ( .x(eop), .a(ncla), .b(csela), .c(asela), .d(i[4]) );
    inv_1 \U891/U1126/U3  ( .x(\U891/reset ), .a(nbReset) );
    inv_1 \U891/U1139/U3  ( .x(\U891/neopack ), .a(eop) );
    nand3_1 \U891/U1131/U9  ( .x(\U891/iay ), .a(\U891/neopack ), .b(
        \U891/naack[0] ), .c(\U891/naack[1] ) );
    nor3_1 \U891/U1128/U27  ( .x(\U891/U1128/nb ), .a(\U891/reset ), .b(\b[3] 
        ), .c(\b[2] ) );
    nor2_1 \U891/U1128/U26  ( .x(\U891/U1128/na ), .a(\b[1] ), .b(\b[0] ) );
    nand2_2 \U891/U1128/U29  ( .x(\U891/ackb ), .a(\U891/U1128/nb ), .b(
        \U891/U1128/na ) );
    nor2_1 \U891/U1133/U5  ( .x(\U891/naack[0] ), .a(\a[3] ), .b(\a[2] ) );
    nor2_1 \U891/U1108/U5  ( .x(\U891/nack ), .a(\U891/acka ), .b(\U891/ackb )
         );
    nor2_1 \U891/U1134/U5  ( .x(\U891/naack[1] ), .a(\a[1] ), .b(\a[0] ) );
    nor2_2 \U891/U914/U6  ( .x(nia), .a(\U891/iay ), .b(\U891/ackb ) );
    nand2_1 \U891/U1130/U5  ( .x(\U891/acka ), .a(\U891/naack[0] ), .b(
        \U891/naack[1] ) );
    ao222_4 \U891/U1121/U1/U1  ( .x(bsela), .a(\U891/nack ), .b(bsel), .c(
        \U891/nack ), .d(bsela), .e(bsel), .f(bsela) );
    ao222_4 \U891/U1120/U1/U1  ( .x(asela), .a(asel), .b(\U891/nack ), .c(asel
        ), .d(asela), .e(\U891/nack ), .f(asela) );
    nor3_1 \U891/U1118_0_/Unr  ( .x(\U891/U1118_0_/nr ), .a(i[0]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_0_/Und  ( .x(\U891/U1118_0_/nd ), .a(i[0]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_0_/U1  ( .x(\U891/U1118_0_/n2 ), .a(\U891/U1118_0_/n2 ), 
        .b(\U891/U1118_0_/nr ), .c(\U891/U1118_0_/nd ) );
    inv_2 \U891/U1118_0_/U3  ( .x(\a[0] ), .a(\U891/U1118_0_/n2 ) );
    nor3_1 \U891/U1118_1_/Unr  ( .x(\U891/U1118_1_/nr ), .a(i[1]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_1_/Und  ( .x(\U891/U1118_1_/nd ), .a(i[1]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_1_/U1  ( .x(\U891/U1118_1_/n2 ), .a(\U891/U1118_1_/n2 ), 
        .b(\U891/U1118_1_/nr ), .c(\U891/U1118_1_/nd ) );
    inv_2 \U891/U1118_1_/U3  ( .x(\a[1] ), .a(\U891/U1118_1_/n2 ) );
    nor3_1 \U891/U1118_2_/Unr  ( .x(\U891/U1118_2_/nr ), .a(i[2]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_2_/Und  ( .x(\U891/U1118_2_/nd ), .a(i[2]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_2_/U1  ( .x(\U891/U1118_2_/n2 ), .a(\U891/U1118_2_/n2 ), 
        .b(\U891/U1118_2_/nr ), .c(\U891/U1118_2_/nd ) );
    inv_2 \U891/U1118_2_/U3  ( .x(\a[2] ), .a(\U891/U1118_2_/n2 ) );
    nor3_1 \U891/U1118_3_/Unr  ( .x(\U891/U1118_3_/nr ), .a(i[3]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_3_/Und  ( .x(\U891/U1118_3_/nd ), .a(i[3]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_3_/U1  ( .x(\U891/U1118_3_/n2 ), .a(\U891/U1118_3_/n2 ), 
        .b(\U891/U1118_3_/nr ), .c(\U891/U1118_3_/nd ) );
    inv_2 \U891/U1118_3_/U3  ( .x(\a[3] ), .a(\U891/U1118_3_/n2 ) );
    nor3_1 \U891/U1117_0_/Unr  ( .x(\U891/U1117_0_/nr ), .a(i[0]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_0_/Und  ( .x(\U891/U1117_0_/nd ), .a(i[0]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_0_/U1  ( .x(\U891/U1117_0_/n2 ), .a(\U891/U1117_0_/n2 ), 
        .b(\U891/U1117_0_/nr ), .c(\U891/U1117_0_/nd ) );
    inv_2 \U891/U1117_0_/U3  ( .x(\b[0] ), .a(\U891/U1117_0_/n2 ) );
    nor3_1 \U891/U1117_1_/Unr  ( .x(\U891/U1117_1_/nr ), .a(i[1]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_1_/Und  ( .x(\U891/U1117_1_/nd ), .a(i[1]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_1_/U1  ( .x(\U891/U1117_1_/n2 ), .a(\U891/U1117_1_/n2 ), 
        .b(\U891/U1117_1_/nr ), .c(\U891/U1117_1_/nd ) );
    inv_2 \U891/U1117_1_/U3  ( .x(\b[1] ), .a(\U891/U1117_1_/n2 ) );
    nor3_1 \U891/U1117_2_/Unr  ( .x(\U891/U1117_2_/nr ), .a(i[2]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_2_/Und  ( .x(\U891/U1117_2_/nd ), .a(i[2]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_2_/U1  ( .x(\U891/U1117_2_/n2 ), .a(\U891/U1117_2_/n2 ), 
        .b(\U891/U1117_2_/nr ), .c(\U891/U1117_2_/nd ) );
    inv_2 \U891/U1117_2_/U3  ( .x(\b[2] ), .a(\U891/U1117_2_/n2 ) );
    nor3_1 \U891/U1117_3_/Unr  ( .x(\U891/U1117_3_/nr ), .a(i[3]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_3_/Und  ( .x(\U891/U1117_3_/nd ), .a(i[3]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_3_/U1  ( .x(\U891/U1117_3_/n2 ), .a(\U891/U1117_3_/n2 ), 
        .b(\U891/U1117_3_/nr ), .c(\U891/U1117_3_/nd ) );
    inv_2 \U891/U1117_3_/U3  ( .x(\b[3] ), .a(\U891/U1117_3_/n2 ) );
    inv_1 \U886/U1126/U3  ( .x(\U886/reset ), .a(nbReset) );
    nor3_1 \U886/U1128/U27  ( .x(\U886/U1128/nb ), .a(\U886/reset ), .b(\f[3] 
        ), .c(\f[2] ) );
    nor2_1 \U886/U1128/U26  ( .x(\U886/U1128/na ), .a(\f[1] ), .b(\f[0] ) );
    nand2_2 \U886/U1128/U29  ( .x(\U886/ackb ), .a(\U886/U1128/nb ), .b(
        \U886/U1128/na ) );
    nor2_1 \U886/U1108/U5  ( .x(\U886/nack ), .a(\U886/acka ), .b(\U886/ackb )
         );
    nor2_2 \U886/U914/U6  ( .x(nba), .a(\U886/acka ), .b(\U886/ackb ) );
    and4_1 \U886/U1127/U25  ( .x(\U886/U1127/n5 ), .a(\U886/U1127/n1 ), .b(
        \U886/U1127/n2 ), .c(\U886/U1127/n3 ), .d(\U886/U1127/n4 ) );
    inv_1 \U886/U1127/U1  ( .x(\U886/U1127/n1 ), .a(\e[3] ) );
    inv_1 \U886/U1127/U2  ( .x(\U886/U1127/n2 ), .a(\e[2] ) );
    inv_1 \U886/U1127/U3  ( .x(\U886/U1127/n3 ), .a(\e[1] ) );
    inv_1 \U886/U1127/U4  ( .x(\U886/U1127/n4 ), .a(\e[0] ) );
    inv_2 \U886/U1127/U5  ( .x(\U886/acka ), .a(\U886/U1127/n5 ) );
    ao222_2 \U886/U1121/U19/U1/U1  ( .x(fsela), .a(\U886/nack ), .b(fsel), .c(
        \U886/nack ), .d(fsela), .e(fsel), .f(fsela) );
    ao222_2 \U886/U1120/U19/U1/U1  ( .x(esela), .a(esel), .b(\U886/nack ), .c(
        esel), .d(esela), .e(\U886/nack ), .f(esela) );
    nor3_1 \U886/U1118_0_/Unr  ( .x(\U886/U1118_0_/nr ), .a(\b[0] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_0_/Und  ( .x(\U886/U1118_0_/nd ), .a(\b[0] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_0_/U1  ( .x(\U886/U1118_0_/n2 ), .a(\U886/U1118_0_/n2 ), 
        .b(\U886/U1118_0_/nr ), .c(\U886/U1118_0_/nd ) );
    inv_2 \U886/U1118_0_/U3  ( .x(\e[0] ), .a(\U886/U1118_0_/n2 ) );
    nor3_1 \U886/U1118_1_/Unr  ( .x(\U886/U1118_1_/nr ), .a(\b[1] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_1_/Und  ( .x(\U886/U1118_1_/nd ), .a(\b[1] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_1_/U1  ( .x(\U886/U1118_1_/n2 ), .a(\U886/U1118_1_/n2 ), 
        .b(\U886/U1118_1_/nr ), .c(\U886/U1118_1_/nd ) );
    inv_2 \U886/U1118_1_/U3  ( .x(\e[1] ), .a(\U886/U1118_1_/n2 ) );
    nor3_1 \U886/U1118_2_/Unr  ( .x(\U886/U1118_2_/nr ), .a(\b[2] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_2_/Und  ( .x(\U886/U1118_2_/nd ), .a(\b[2] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_2_/U1  ( .x(\U886/U1118_2_/n2 ), .a(\U886/U1118_2_/n2 ), 
        .b(\U886/U1118_2_/nr ), .c(\U886/U1118_2_/nd ) );
    inv_2 \U886/U1118_2_/U3  ( .x(\e[2] ), .a(\U886/U1118_2_/n2 ) );
    nor3_1 \U886/U1118_3_/Unr  ( .x(\U886/U1118_3_/nr ), .a(\b[3] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_3_/Und  ( .x(\U886/U1118_3_/nd ), .a(\b[3] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_3_/U1  ( .x(\U886/U1118_3_/n2 ), .a(\U886/U1118_3_/n2 ), 
        .b(\U886/U1118_3_/nr ), .c(\U886/U1118_3_/nd ) );
    inv_2 \U886/U1118_3_/U3  ( .x(\e[3] ), .a(\U886/U1118_3_/n2 ) );
    nor3_1 \U886/U1117_0_/Unr  ( .x(\U886/U1117_0_/nr ), .a(\b[0] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_0_/Und  ( .x(\U886/U1117_0_/nd ), .a(\b[0] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_0_/U1  ( .x(\U886/U1117_0_/n2 ), .a(\U886/U1117_0_/n2 ), 
        .b(\U886/U1117_0_/nr ), .c(\U886/U1117_0_/nd ) );
    inv_2 \U886/U1117_0_/U3  ( .x(\f[0] ), .a(\U886/U1117_0_/n2 ) );
    nor3_1 \U886/U1117_1_/Unr  ( .x(\U886/U1117_1_/nr ), .a(\b[1] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_1_/Und  ( .x(\U886/U1117_1_/nd ), .a(\b[1] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_1_/U1  ( .x(\U886/U1117_1_/n2 ), .a(\U886/U1117_1_/n2 ), 
        .b(\U886/U1117_1_/nr ), .c(\U886/U1117_1_/nd ) );
    inv_2 \U886/U1117_1_/U3  ( .x(\f[1] ), .a(\U886/U1117_1_/n2 ) );
    nor3_1 \U886/U1117_2_/Unr  ( .x(\U886/U1117_2_/nr ), .a(\b[2] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_2_/Und  ( .x(\U886/U1117_2_/nd ), .a(\b[2] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_2_/U1  ( .x(\U886/U1117_2_/n2 ), .a(\U886/U1117_2_/n2 ), 
        .b(\U886/U1117_2_/nr ), .c(\U886/U1117_2_/nd ) );
    inv_2 \U886/U1117_2_/U3  ( .x(\f[2] ), .a(\U886/U1117_2_/n2 ) );
    nor3_1 \U886/U1117_3_/Unr  ( .x(\U886/U1117_3_/nr ), .a(\b[3] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_3_/Und  ( .x(\U886/U1117_3_/nd ), .a(\b[3] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_3_/U1  ( .x(\U886/U1117_3_/n2 ), .a(\U886/U1117_3_/n2 ), 
        .b(\U886/U1117_3_/nr ), .c(\U886/U1117_3_/nd ) );
    inv_2 \U886/U1117_3_/U3  ( .x(\f[3] ), .a(\U886/U1117_3_/n2 ) );
    inv_1 \U884/U1126/U3  ( .x(\U884/reset ), .a(nbReset) );
    nor3_1 \U884/U1128/U27  ( .x(\U884/U1128/nb ), .a(\U884/reset ), .b(\d[3] 
        ), .c(\d[2] ) );
    nor2_1 \U884/U1128/U26  ( .x(\U884/U1128/na ), .a(\d[1] ), .b(\d[0] ) );
    nand2_2 \U884/U1128/U29  ( .x(\U884/ackb ), .a(\U884/U1128/nb ), .b(
        \U884/U1128/na ) );
    nor2_1 \U884/U1108/U5  ( .x(\U884/nack ), .a(\U884/acka ), .b(\U884/ackb )
         );
    nor2_2 \U884/U914/U6  ( .x(naa), .a(\U884/acka ), .b(\U884/ackb ) );
    and4_1 \U884/U1127/U25  ( .x(\U884/U1127/n5 ), .a(\U884/U1127/n1 ), .b(
        \U884/U1127/n2 ), .c(\U884/U1127/n3 ), .d(\U884/U1127/n4 ) );
    inv_1 \U884/U1127/U1  ( .x(\U884/U1127/n1 ), .a(\c[3] ) );
    inv_1 \U884/U1127/U2  ( .x(\U884/U1127/n2 ), .a(\c[2] ) );
    inv_1 \U884/U1127/U3  ( .x(\U884/U1127/n3 ), .a(\c[1] ) );
    inv_1 \U884/U1127/U4  ( .x(\U884/U1127/n4 ), .a(\c[0] ) );
    inv_2 \U884/U1127/U5  ( .x(\U884/acka ), .a(\U884/U1127/n5 ) );
    ao222_2 \U884/U1121/U19/U1/U1  ( .x(dsela), .a(\U884/nack ), .b(dsel), .c(
        \U884/nack ), .d(dsela), .e(dsel), .f(dsela) );
    ao222_2 \U884/U1120/U19/U1/U1  ( .x(csela), .a(csel), .b(\U884/nack ), .c(
        csel), .d(csela), .e(\U884/nack ), .f(csela) );
    nor3_1 \U884/U1118_0_/Unr  ( .x(\U884/U1118_0_/nr ), .a(\a[0] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_0_/Und  ( .x(\U884/U1118_0_/nd ), .a(\a[0] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_0_/U1  ( .x(\U884/U1118_0_/n2 ), .a(\U884/U1118_0_/n2 ), 
        .b(\U884/U1118_0_/nr ), .c(\U884/U1118_0_/nd ) );
    inv_2 \U884/U1118_0_/U3  ( .x(\c[0] ), .a(\U884/U1118_0_/n2 ) );
    nor3_1 \U884/U1118_1_/Unr  ( .x(\U884/U1118_1_/nr ), .a(\a[1] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_1_/Und  ( .x(\U884/U1118_1_/nd ), .a(\a[1] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_1_/U1  ( .x(\U884/U1118_1_/n2 ), .a(\U884/U1118_1_/n2 ), 
        .b(\U884/U1118_1_/nr ), .c(\U884/U1118_1_/nd ) );
    inv_2 \U884/U1118_1_/U3  ( .x(\c[1] ), .a(\U884/U1118_1_/n2 ) );
    nor3_1 \U884/U1118_2_/Unr  ( .x(\U884/U1118_2_/nr ), .a(\a[2] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_2_/Und  ( .x(\U884/U1118_2_/nd ), .a(\a[2] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_2_/U1  ( .x(\U884/U1118_2_/n2 ), .a(\U884/U1118_2_/n2 ), 
        .b(\U884/U1118_2_/nr ), .c(\U884/U1118_2_/nd ) );
    inv_2 \U884/U1118_2_/U3  ( .x(\c[2] ), .a(\U884/U1118_2_/n2 ) );
    nor3_1 \U884/U1118_3_/Unr  ( .x(\U884/U1118_3_/nr ), .a(\a[3] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_3_/Und  ( .x(\U884/U1118_3_/nd ), .a(\a[3] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_3_/U1  ( .x(\U884/U1118_3_/n2 ), .a(\U884/U1118_3_/n2 ), 
        .b(\U884/U1118_3_/nr ), .c(\U884/U1118_3_/nd ) );
    inv_2 \U884/U1118_3_/U3  ( .x(\c[3] ), .a(\U884/U1118_3_/n2 ) );
    nor3_1 \U884/U1117_0_/Unr  ( .x(\U884/U1117_0_/nr ), .a(\a[0] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_0_/Und  ( .x(\U884/U1117_0_/nd ), .a(\a[0] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_0_/U1  ( .x(\U884/U1117_0_/n2 ), .a(\U884/U1117_0_/n2 ), 
        .b(\U884/U1117_0_/nr ), .c(\U884/U1117_0_/nd ) );
    inv_2 \U884/U1117_0_/U3  ( .x(\d[0] ), .a(\U884/U1117_0_/n2 ) );
    nor3_1 \U884/U1117_1_/Unr  ( .x(\U884/U1117_1_/nr ), .a(\a[1] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_1_/Und  ( .x(\U884/U1117_1_/nd ), .a(\a[1] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_1_/U1  ( .x(\U884/U1117_1_/n2 ), .a(\U884/U1117_1_/n2 ), 
        .b(\U884/U1117_1_/nr ), .c(\U884/U1117_1_/nd ) );
    inv_2 \U884/U1117_1_/U3  ( .x(\d[1] ), .a(\U884/U1117_1_/n2 ) );
    nor3_1 \U884/U1117_2_/Unr  ( .x(\U884/U1117_2_/nr ), .a(\a[2] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_2_/Und  ( .x(\U884/U1117_2_/nd ), .a(\a[2] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_2_/U1  ( .x(\U884/U1117_2_/n2 ), .a(\U884/U1117_2_/n2 ), 
        .b(\U884/U1117_2_/nr ), .c(\U884/U1117_2_/nd ) );
    inv_2 \U884/U1117_2_/U3  ( .x(\d[2] ), .a(\U884/U1117_2_/n2 ) );
    nor3_1 \U884/U1117_3_/Unr  ( .x(\U884/U1117_3_/nr ), .a(\a[3] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_3_/Und  ( .x(\U884/U1117_3_/nd ), .a(\a[3] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_3_/U1  ( .x(\U884/U1117_3_/n2 ), .a(\U884/U1117_3_/n2 ), 
        .b(\U884/U1117_3_/nr ), .c(\U884/U1117_3_/nd ) );
    inv_2 \U884/U1117_3_/U3  ( .x(\d[3] ), .a(\U884/U1117_3_/n2 ) );
    nand2_1 \U888/U1128/U5  ( .x(\U888/s ), .a(\U888/r ), .b(\U888/nback ) );
    nand2_1 \U888/U1103/U5  ( .x(\U888/r ), .a(\U888/naack ), .b(\U888/s ) );
    inv_1 \U888/U1111/U3  ( .x(\U888/reset ), .a(nbReset) );
    inv_1 \U888/U1112/U3  ( .x(\U888/naack ), .a(esela) );
    nor2_1 \U888/U1127/U5  ( .x(\U888/nback ), .a(fsela), .b(\U888/reset ) );
    and2_2 \U888/U1129/U8  ( .x(esel), .a(\U888/nback ), .b(\U888/s ) );
    and2_2 \U888/U1124/U8  ( .x(fsel), .a(\U888/r ), .b(\U888/naack ) );
    nand2_1 \U887/U1128/U5  ( .x(\U887/s ), .a(\U887/r ), .b(\U887/nback ) );
    nand2_1 \U887/U1103/U5  ( .x(\U887/r ), .a(\U887/naack ), .b(\U887/s ) );
    inv_1 \U887/U1111/U3  ( .x(\U887/reset ), .a(nbReset) );
    inv_1 \U887/U1112/U3  ( .x(\U887/naack ), .a(csela) );
    nor2_1 \U887/U1127/U5  ( .x(\U887/nback ), .a(dsela), .b(\U887/reset ) );
    and2_2 \U887/U1129/U8  ( .x(csel), .a(\U887/nback ), .b(\U887/s ) );
    and2_2 \U887/U1124/U8  ( .x(dsel), .a(\U887/r ), .b(\U887/naack ) );
    nand2_1 \U885/U1128/U5  ( .x(\U885/s ), .a(\U885/r ), .b(\U885/nback ) );
    nand2_1 \U885/U1103/U5  ( .x(\U885/r ), .a(\U885/naack ), .b(\U885/s ) );
    inv_1 \U885/U1111/U3  ( .x(\U885/reset ), .a(nbReset) );
    inv_1 \U885/U1112/U3  ( .x(\U885/naack ), .a(asela) );
    nor2_1 \U885/U1127/U5  ( .x(\U885/nback ), .a(bsela), .b(\U885/reset ) );
    and2_2 \U885/U1129/U8  ( .x(asel), .a(\U885/nback ), .b(\U885/s ) );
    and2_2 \U885/U1124/U8  ( .x(bsel), .a(\U885/r ), .b(\U885/naack ) );
    nor3_1 \U877/U594/U7  ( .x(\U877/x ), .a(ol[7]), .b(\U877/reset ), .c(oh
        [7]) );
    nor3_1 \U877/U593/U7  ( .x(\U877/y ), .a(ol[6]), .b(\U877/reset ), .c(oh
        [6]) );
    inv_1 \U877/U604/U3  ( .x(\U877/reset ), .a(nbReset) );
    oa31_1 \U877/U590/U25/U1/Uclr  ( .x(\U877/U590/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[1] ), .d(oh[6]) );
    oaoi211_1 \U877/U590/U25/U1/Uaoi  ( .x(\U877/U590/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[1] ), .c(n1), .d(\U877/U590/U25/U1/clr ) );
    inv_2 \U877/U590/U25/U1/Ui  ( .x(oh[6]), .a(\U877/U590/U25/U1/ob ) );
    oa31_1 \U877/U589/U25/U1/Uclr  ( .x(\U877/U589/U25/U1/clr ), .a(net135), 
        .b(\cl[1] ), .c(\cl[0] ), .d(ol[7]) );
    oaoi211_1 \U877/U589/U25/U1/Uaoi  ( .x(\U877/U589/U25/U1/ob ), .a(\cl[1] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U589/U25/U1/clr ) );
    inv_2 \U877/U589/U25/U1/Ui  ( .x(ol[7]), .a(\U877/U589/U25/U1/ob ) );
    oa31_1 \U877/U588/U25/U1/Uclr  ( .x(\U877/U588/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[2] ), .d(oh[7]) );
    oaoi211_1 \U877/U588/U25/U1/Uaoi  ( .x(\U877/U588/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[2] ), .c(n1), .d(\U877/U588/U25/U1/clr ) );
    inv_2 \U877/U588/U25/U1/Ui  ( .x(oh[7]), .a(\U877/U588/U25/U1/ob ) );
    oa31_1 \U877/U591/U25/U1/Uclr  ( .x(\U877/U591/U25/U1/clr ), .a(net135), 
        .b(\cl[2] ), .c(\cl[0] ), .d(ol[6]) );
    oaoi211_1 \U877/U591/U25/U1/Uaoi  ( .x(\U877/U591/U25/U1/ob ), .a(\cl[2] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U591/U25/U1/clr ) );
    inv_2 \U877/U591/U25/U1/Ui  ( .x(ol[6]), .a(\U877/U591/U25/U1/ob ) );
    ao222_2 \U877/U592/U19/U1/U1  ( .x(ncla), .a(\U877/x ), .b(\U877/y ), .c(
        \U877/x ), .d(ncla), .e(\U877/y ), .f(ncla) );
    nor3_1 \U876/U594/U7  ( .x(\U876/x ), .a(ol[3]), .b(\U876/reset ), .c(oh
        [3]) );
    nor3_1 \U876/U593/U7  ( .x(\U876/y ), .a(ol[2]), .b(\U876/reset ), .c(oh
        [2]) );
    inv_1 \U876/U604/U3  ( .x(\U876/reset ), .a(nbReset) );
    oa31_1 \U876/U590/U25/U1/Uclr  ( .x(\U876/U590/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[1] ), .d(oh[2]) );
    oaoi211_1 \U876/U590/U25/U1/Uaoi  ( .x(\U876/U590/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[1] ), .c(n1), .d(\U876/U590/U25/U1/clr ) );
    inv_2 \U876/U590/U25/U1/Ui  ( .x(oh[2]), .a(\U876/U590/U25/U1/ob ) );
    oa31_1 \U876/U589/U25/U1/Uclr  ( .x(\U876/U589/U25/U1/clr ), .a(net135), 
        .b(\d[1] ), .c(\d[0] ), .d(ol[3]) );
    oaoi211_1 \U876/U589/U25/U1/Uaoi  ( .x(\U876/U589/U25/U1/ob ), .a(\d[1] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U589/U25/U1/clr ) );
    inv_2 \U876/U589/U25/U1/Ui  ( .x(ol[3]), .a(\U876/U589/U25/U1/ob ) );
    oa31_1 \U876/U588/U25/U1/Uclr  ( .x(\U876/U588/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[2] ), .d(oh[3]) );
    oaoi211_1 \U876/U588/U25/U1/Uaoi  ( .x(\U876/U588/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[2] ), .c(n1), .d(\U876/U588/U25/U1/clr ) );
    inv_2 \U876/U588/U25/U1/Ui  ( .x(oh[3]), .a(\U876/U588/U25/U1/ob ) );
    oa31_1 \U876/U591/U25/U1/Uclr  ( .x(\U876/U591/U25/U1/clr ), .a(net135), 
        .b(\d[2] ), .c(\d[0] ), .d(ol[2]) );
    oaoi211_1 \U876/U591/U25/U1/Uaoi  ( .x(\U876/U591/U25/U1/ob ), .a(\d[2] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U591/U25/U1/clr ) );
    inv_2 \U876/U591/U25/U1/Ui  ( .x(ol[2]), .a(\U876/U591/U25/U1/ob ) );
    ao222_2 \U876/U592/U19/U1/U1  ( .x(nda), .a(\U876/x ), .b(\U876/y ), .c(
        \U876/x ), .d(nda), .e(\U876/y ), .f(nda) );
    nor3_1 \U2/U594/U7  ( .x(\U2/x ), .a(ol[1]), .b(\U2/reset ), .c(oh[1]) );
    nor3_1 \U2/U593/U7  ( .x(\U2/y ), .a(ol[0]), .b(\U2/reset ), .c(oh[0]) );
    inv_1 \U2/U604/U3  ( .x(\U2/reset ), .a(nbReset) );
    oa31_1 \U2/U590/U25/U1/Uclr  ( .x(\U2/U590/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[1] ), .d(oh[0]) );
    oaoi211_1 \U2/U590/U25/U1/Uaoi  ( .x(\U2/U590/U25/U1/ob ), .a(\f[3] ), .b(
        \f[1] ), .c(n1), .d(\U2/U590/U25/U1/clr ) );
    inv_2 \U2/U590/U25/U1/Ui  ( .x(oh[0]), .a(\U2/U590/U25/U1/ob ) );
    oa31_1 \U2/U589/U25/U1/Uclr  ( .x(\U2/U589/U25/U1/clr ), .a(net135), .b(
        \f[1] ), .c(\f[0] ), .d(ol[1]) );
    oaoi211_1 \U2/U589/U25/U1/Uaoi  ( .x(\U2/U589/U25/U1/ob ), .a(\f[1] ), .b(
        \f[0] ), .c(n1), .d(\U2/U589/U25/U1/clr ) );
    inv_2 \U2/U589/U25/U1/Ui  ( .x(ol[1]), .a(\U2/U589/U25/U1/ob ) );
    oa31_1 \U2/U588/U25/U1/Uclr  ( .x(\U2/U588/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[2] ), .d(oh[1]) );
    oaoi211_1 \U2/U588/U25/U1/Uaoi  ( .x(\U2/U588/U25/U1/ob ), .a(\f[3] ), .b(
        \f[2] ), .c(n1), .d(\U2/U588/U25/U1/clr ) );
    inv_2 \U2/U588/U25/U1/Ui  ( .x(oh[1]), .a(\U2/U588/U25/U1/ob ) );
    oa31_1 \U2/U591/U25/U1/Uclr  ( .x(\U2/U591/U25/U1/clr ), .a(net135), .b(
        \f[2] ), .c(\f[0] ), .d(ol[0]) );
    oaoi211_1 \U2/U591/U25/U1/Uaoi  ( .x(\U2/U591/U25/U1/ob ), .a(\f[2] ), .b(
        \f[0] ), .c(n1), .d(\U2/U591/U25/U1/clr ) );
    inv_2 \U2/U591/U25/U1/Ui  ( .x(ol[0]), .a(\U2/U591/U25/U1/ob ) );
    ao222_2 \U2/U592/U19/U1/U1  ( .x(nfa), .a(\U2/x ), .b(\U2/y ), .c(\U2/x ), 
        .d(nfa), .e(\U2/y ), .f(nfa) );
    nor3_1 \U1/U594/U7  ( .x(\U1/x ), .a(ol[5]), .b(\U1/reset ), .c(oh[5]) );
    nor3_1 \U1/U593/U7  ( .x(\U1/y ), .a(ol[4]), .b(\U1/reset ), .c(oh[4]) );
    inv_1 \U1/U604/U3  ( .x(\U1/reset ), .a(nbReset) );
    oa31_1 \U1/U590/U25/U1/Uclr  ( .x(\U1/U590/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[1] ), .d(oh[4]) );
    oaoi211_1 \U1/U590/U25/U1/Uaoi  ( .x(\U1/U590/U25/U1/ob ), .a(\e[3] ), .b(
        \e[1] ), .c(n1), .d(\U1/U590/U25/U1/clr ) );
    inv_2 \U1/U590/U25/U1/Ui  ( .x(oh[4]), .a(\U1/U590/U25/U1/ob ) );
    oa31_1 \U1/U589/U25/U1/Uclr  ( .x(\U1/U589/U25/U1/clr ), .a(net135), .b(
        \e[1] ), .c(\e[0] ), .d(ol[5]) );
    oaoi211_1 \U1/U589/U25/U1/Uaoi  ( .x(\U1/U589/U25/U1/ob ), .a(\e[1] ), .b(
        \e[0] ), .c(n1), .d(\U1/U589/U25/U1/clr ) );
    inv_2 \U1/U589/U25/U1/Ui  ( .x(ol[5]), .a(\U1/U589/U25/U1/ob ) );
    oa31_1 \U1/U588/U25/U1/Uclr  ( .x(\U1/U588/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[2] ), .d(oh[5]) );
    oaoi211_1 \U1/U588/U25/U1/Uaoi  ( .x(\U1/U588/U25/U1/ob ), .a(\e[3] ), .b(
        \e[2] ), .c(n1), .d(\U1/U588/U25/U1/clr ) );
    inv_2 \U1/U588/U25/U1/Ui  ( .x(oh[5]), .a(\U1/U588/U25/U1/ob ) );
    oa31_1 \U1/U591/U25/U1/Uclr  ( .x(\U1/U591/U25/U1/clr ), .a(net135), .b(
        \e[2] ), .c(\e[0] ), .d(ol[4]) );
    oaoi211_1 \U1/U591/U25/U1/Uaoi  ( .x(\U1/U591/U25/U1/ob ), .a(\e[2] ), .b(
        \e[0] ), .c(n1), .d(\U1/U591/U25/U1/clr ) );
    inv_2 \U1/U591/U25/U1/Ui  ( .x(ol[4]), .a(\U1/U591/U25/U1/ob ) );
    ao222_2 \U1/U592/U19/U1/U1  ( .x(nea), .a(\U1/x ), .b(\U1/y ), .c(\U1/x ), 
        .d(nea), .e(\U1/y ), .f(nea) );
    and3_4 \U881/U20/U9  ( .x(nca), .a(\U881/nack[1] ), .b(\U881/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U881/U18/U5  ( .x(\U881/nack[0] ), .a(\cl[3] ), .b(\cl[0] ) );
    nor2_1 \U881/U19/U5  ( .x(\U881/nack[1] ), .a(\cl[1] ), .b(\cl[2] ) );
    ao222_2 \U881/U15_0_/U19/U1/U1  ( .x(\cl[0] ), .a(\c[0] ), .b(ncla), .c(
        \c[0] ), .d(\cl[0] ), .e(ncla), .f(\cl[0] ) );
    ao222_2 \U881/U15_1_/U19/U1/U1  ( .x(\cl[1] ), .a(\c[1] ), .b(ncla), .c(
        \c[1] ), .d(\cl[1] ), .e(ncla), .f(\cl[1] ) );
    ao222_2 \U881/U15_2_/U19/U1/U1  ( .x(\cl[2] ), .a(\c[2] ), .b(ncla), .c(
        \c[2] ), .d(\cl[2] ), .e(ncla), .f(\cl[2] ) );
    ao222_2 \U881/U15_3_/U19/U1/U1  ( .x(\cl[3] ), .a(\c[3] ), .b(ncla), .c(
        \c[3] ), .d(\cl[3] ), .e(ncla), .f(\cl[3] ) );
    and2_5 U1 ( .x(n1), .a(nbReset), .b(noa) );
    and2_3 U2 ( .x(net135), .a(nbReset), .b(noa) );
endmodule


module chain_dr2fr_byte_4 ( eop_ack, ia, o, eop, ih, il, nReset, noa );
output [4:0] o;
input  [7:0] ih;
input  [7:0] il;
input  eop, nReset, noa;
output eop_ack, ia;
    wire eop_pass, nhighack, nlowack, \twobitack[2] , \twobitack[3] , 
        \twobitack[0] , \twobitack[1] , xsel, ysel, nxa, nyla, nbReset, nya, 
        \y[3] , \y[2] , \y[1] , \y[0] , \yl[3] , \yl[2] , \yl[1] , \yl[0] , 
        \cdh[0] , \cdh[1] , \cdl[0] , \cdl[1] , net193, \cdh[2] , \cdh[3] , 
        \cdl[2] , \cdl[3] , net195, bsel, dsel, nba, bg, nda, dg, asel, csel, 
        naa, ag, nca, cg, \d[3] , \d[2] , \d[1] , \d[0] , \b[3] , \b[2] , 
        \b[1] , \b[0] , \x[3] , \x[2] , \x[1] , \x[0] , \c[3] , \c[2] , \c[1] , 
        \c[0] , \a[3] , \a[2] , \a[1] , \a[0] , net194, net199, \U1018/Z , 
        \U1270/net190 , \U1270/net191 , \U1270/net192 , \U1270/net189 , 
        \U1270/U1141/Z , \U1268/net190 , \U1268/net191 , \U1268/net192 , 
        \U1268/net189 , \U1268/U1141/Z , \U1224/nack[0] , \U1224/nack[1] , 
        \U1224/net4 , \U1224/U1125/U28/U1/clr , \U1224/U1125/U28/U1/set , 
        \U1224/U1122/U28/U1/clr , \U1224/U1122/U28/U1/set , 
        \U1224/U916_0_/U25/U1/clr , \U1224/U916_0_/U25/U1/ob , 
        \U1224/U916_1_/U25/U1/clr , \U1224/U916_1_/U25/U1/ob , 
        \U1224/U916_2_/U25/U1/clr , \U1224/U916_2_/U25/U1/ob , 
        \U1224/U916_3_/U25/U1/clr , \U1224/U916_3_/U25/U1/ob , \U1209/nack[0] , 
        \U1209/nack[1] , \U1209/net4 , \U1209/U1125/U28/U1/clr , 
        \U1209/U1125/U28/U1/set , \U1209/U1122/U28/U1/clr , 
        \U1209/U1122/U28/U1/set , \U1209/U916_0_/U25/U1/clr , 
        \U1209/U916_0_/U25/U1/ob , \U1209/U916_1_/U25/U1/clr , 
        \U1209/U916_1_/U25/U1/ob , \U1209/U916_2_/U25/U1/clr , 
        \U1209/U916_2_/U25/U1/ob , \U1209/U916_3_/U25/U1/clr , 
        \U1209/U916_3_/U25/U1/ob , \U1213/nack[0] , \U1213/nack[1] , 
        \U1213/net4 , \U1213/U1125/U28/U1/clr , \U1213/U1125/U28/U1/set , 
        \U1213/U1122/U28/U1/clr , \U1213/U1122/U28/U1/set , 
        \U1213/U916_0_/U25/U1/clr , \U1213/U916_0_/U25/U1/ob , 
        \U1213/U916_1_/U25/U1/clr , \U1213/U916_1_/U25/U1/ob , 
        \U1213/U916_2_/U25/U1/clr , \U1213/U916_2_/U25/U1/ob , 
        \U1213/U916_3_/U25/U1/clr , \U1213/U916_3_/U25/U1/ob , \U1296/ng , 
        \U1296/U1384/Z , \U1296/U1386/U25/U1/clr , \U1296/U1386/U25/U1/ob , 
        \U1298/ng , \U1298/U1384/Z , \U1298/U1386/U25/U1/clr , 
        \U1298/U1386/U25/U1/ob , \U1306/ng , \U1306/U1384/Z , 
        \U1306/U1386/U25/U1/clr , \U1306/U1386/U25/U1/ob , \U1295/ng , 
        \U1295/U1384/Z , \U1295/U1386/U25/U1/clr , \U1295/U1386/U25/U1/ob , 
        \U1297/s , \U1297/nback , \U1297/r , \U1297/naack , \U1297/reset , 
        \U1297/U1128/U28/U1/clr , \U1297/U1128/U28/U1/set , 
        \U1297/U1127/U28/U1/clr , \U1297/U1127/U28/U1/set , \U1300/s , 
        \U1300/nback , \U1300/r , \U1300/naack , \U1300/reset , 
        \U1300/U1128/U28/U1/clr , \U1300/U1128/U28/U1/set , 
        \U1300/U1127/U28/U1/clr , \U1300/U1127/U28/U1/set , \U1289/bnreset , 
        \U1289/U1150/U28/U1/clr , \U1289/U1150/U28/U1/set , 
        \U1289/U1152/U28/U1/clr , \U1289/U1152/U28/U1/set , 
        \U1289/U1149/U28/U1/clr , \U1289/U1149/U28/U1/set , 
        \U1289/U1151/U28/U1/clr , \U1289/U1151/U28/U1/set , 
        \U1289/U1148/net190 , \U1289/U1148/net191 , \U1289/U1148/net192 , 
        \U1289/U1148/net189 , \U1289/U1148/U1141/Z , \U1271/bnreset , 
        \U1271/U1150/U28/U1/clr , \U1271/U1150/U28/U1/set , 
        \U1271/U1152/U28/U1/clr , \U1271/U1152/U28/U1/set , 
        \U1271/U1149/U28/U1/clr , \U1271/U1149/U28/U1/set , 
        \U1271/U1151/U28/U1/clr , \U1271/U1151/U28/U1/set , 
        \U1271/U1148/net190 , \U1271/U1148/net191 , \U1271/U1148/net192 , 
        \U1271/U1148/net189 , \U1271/U1148/U1141/Z , \U1225/naack , \U1225/r , 
        \U1225/s , \U1225/nback , \U1225/reset , \U1308/nack[1] , 
        \U1308/nack[0] ;
    assign o[4] = eop_ack;
    buf_2 U1231 ( .x(nbReset), .a(nReset) );
    and3_1 \U1194/U9  ( .x(eop_pass), .a(nxa), .b(naa), .c(eop) );
    ao222_1 \U1301/U18/U1/U1  ( .x(nlowack), .a(\twobitack[0] ), .b(
        \twobitack[1] ), .c(\twobitack[0] ), .d(nlowack), .e(\twobitack[1] ), 
        .f(nlowack) );
    ao222_1 \U1302/U18/U1/U1  ( .x(nhighack), .a(\twobitack[2] ), .b(
        \twobitack[3] ), .c(\twobitack[2] ), .d(nhighack), .e(\twobitack[3] ), 
        .f(nhighack) );
    aoi222_1 \U1018/U30/U1  ( .x(ia), .a(nhighack), .b(nlowack), .c(nhighack), 
        .d(\U1018/Z ), .e(nlowack), .f(\U1018/Z ) );
    inv_1 \U1018/U30/Uinv  ( .x(\U1018/Z ), .a(ia) );
    ao222_2 \U1038/U19/U1/U1  ( .x(eop_ack), .a(eop_pass), .b(noa), .c(
        eop_pass), .d(eop_ack), .e(noa), .f(eop_ack) );
    inv_1 \U1270/U1147/U3  ( .x(\U1270/net189 ), .a(nbReset) );
    nor2_1 \U1270/U582/U5  ( .x(\U1270/net192 ), .a(il[4]), .b(ih[4]) );
    nor2_1 \U1270/U580/U5  ( .x(\U1270/net191 ), .a(il[5]), .b(ih[5]) );
    nor2_2 \U1270/U1146/U6  ( .x(net199), .a(\U1270/net190 ), .b(
        \U1270/net189 ) );
    aoi222_1 \U1270/U1141/U30/U1  ( .x(\U1270/net190 ), .a(\U1270/net191 ), 
        .b(\U1270/net192 ), .c(\U1270/net191 ), .d(\U1270/U1141/Z ), .e(
        \U1270/net192 ), .f(\U1270/U1141/Z ) );
    inv_1 \U1270/U1141/U30/Uinv  ( .x(\U1270/U1141/Z ), .a(\U1270/net190 ) );
    inv_1 \U1268/U1147/U3  ( .x(\U1268/net189 ), .a(nbReset) );
    nor2_1 \U1268/U582/U5  ( .x(\U1268/net192 ), .a(il[6]), .b(ih[6]) );
    nor2_1 \U1268/U580/U5  ( .x(\U1268/net191 ), .a(il[7]), .b(ih[7]) );
    nor2_2 \U1268/U1146/U6  ( .x(net194), .a(\U1268/net190 ), .b(
        \U1268/net189 ) );
    aoi222_1 \U1268/U1141/U30/U1  ( .x(\U1268/net190 ), .a(\U1268/net191 ), 
        .b(\U1268/net192 ), .c(\U1268/net191 ), .d(\U1268/U1141/Z ), .e(
        \U1268/net192 ), .f(\U1268/U1141/Z ) );
    inv_1 \U1268/U1141/U30/Uinv  ( .x(\U1268/U1141/Z ), .a(\U1268/net190 ) );
    nor2_1 \U1224/U1128/U5  ( .x(\U1224/nack[0] ), .a(\x[3] ), .b(\x[2] ) );
    nor3_1 \U1224/U1127/U7  ( .x(\U1224/nack[1] ), .a(\x[1] ), .b(\U1224/net4 
        ), .c(\x[0] ) );
    inv_1 \U1224/U907/U3  ( .x(\U1224/net4 ), .a(nbReset) );
    aoai211_1 \U1224/U1125/U28/U1/U1  ( .x(\U1224/U1125/U28/U1/clr ), .a(
        \U1224/nack[1] ), .b(\U1224/nack[0] ), .c(asel), .d(naa) );
    nand3_1 \U1224/U1125/U28/U1/U2  ( .x(\U1224/U1125/U28/U1/set ), .a(asel), 
        .b(\U1224/nack[1] ), .c(\U1224/nack[0] ) );
    nand2_2 \U1224/U1125/U28/U1/U3  ( .x(naa), .a(\U1224/U1125/U28/U1/clr ), 
        .b(\U1224/U1125/U28/U1/set ) );
    aoai211_1 \U1224/U1122/U28/U1/U1  ( .x(\U1224/U1122/U28/U1/clr ), .a(
        \U1224/nack[0] ), .b(\U1224/nack[1] ), .c(csel), .d(nca) );
    nand3_1 \U1224/U1122/U28/U1/U2  ( .x(\U1224/U1122/U28/U1/set ), .a(csel), 
        .b(\U1224/nack[0] ), .c(\U1224/nack[1] ) );
    nand2_2 \U1224/U1122/U28/U1/U3  ( .x(nca), .a(\U1224/U1122/U28/U1/clr ), 
        .b(\U1224/U1122/U28/U1/set ) );
    oa31_1 \U1224/U916_0_/U25/U1/Uclr  ( .x(\U1224/U916_0_/U25/U1/clr ), .a(
        nxa), .b(\a[0] ), .c(\c[0] ), .d(\x[0] ) );
    oaoi211_1 \U1224/U916_0_/U25/U1/Uaoi  ( .x(\U1224/U916_0_/U25/U1/ob ), .a(
        \a[0] ), .b(\c[0] ), .c(nxa), .d(\U1224/U916_0_/U25/U1/clr ) );
    inv_2 \U1224/U916_0_/U25/U1/Ui  ( .x(\x[0] ), .a(\U1224/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_1_/U25/U1/Uclr  ( .x(\U1224/U916_1_/U25/U1/clr ), .a(
        nxa), .b(\a[1] ), .c(\c[1] ), .d(\x[1] ) );
    oaoi211_1 \U1224/U916_1_/U25/U1/Uaoi  ( .x(\U1224/U916_1_/U25/U1/ob ), .a(
        \a[1] ), .b(\c[1] ), .c(nxa), .d(\U1224/U916_1_/U25/U1/clr ) );
    inv_2 \U1224/U916_1_/U25/U1/Ui  ( .x(\x[1] ), .a(\U1224/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_2_/U25/U1/Uclr  ( .x(\U1224/U916_2_/U25/U1/clr ), .a(
        nxa), .b(\a[2] ), .c(\c[2] ), .d(\x[2] ) );
    oaoi211_1 \U1224/U916_2_/U25/U1/Uaoi  ( .x(\U1224/U916_2_/U25/U1/ob ), .a(
        \a[2] ), .b(\c[2] ), .c(nxa), .d(\U1224/U916_2_/U25/U1/clr ) );
    inv_2 \U1224/U916_2_/U25/U1/Ui  ( .x(\x[2] ), .a(\U1224/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_3_/U25/U1/Uclr  ( .x(\U1224/U916_3_/U25/U1/clr ), .a(
        nxa), .b(\a[3] ), .c(\c[3] ), .d(\x[3] ) );
    oaoi211_1 \U1224/U916_3_/U25/U1/Uaoi  ( .x(\U1224/U916_3_/U25/U1/ob ), .a(
        \a[3] ), .b(\c[3] ), .c(nxa), .d(\U1224/U916_3_/U25/U1/clr ) );
    inv_2 \U1224/U916_3_/U25/U1/Ui  ( .x(\x[3] ), .a(\U1224/U916_3_/U25/U1/ob 
        ) );
    nor2_1 \U1209/U1128/U5  ( .x(\U1209/nack[0] ), .a(o[3]), .b(o[2]) );
    nor3_1 \U1209/U1127/U7  ( .x(\U1209/nack[1] ), .a(o[1]), .b(\U1209/net4 ), 
        .c(o[0]) );
    inv_1 \U1209/U907/U3  ( .x(\U1209/net4 ), .a(nbReset) );
    aoai211_1 \U1209/U1125/U28/U1/U1  ( .x(\U1209/U1125/U28/U1/clr ), .a(
        \U1209/nack[1] ), .b(\U1209/nack[0] ), .c(xsel), .d(nxa) );
    nand3_1 \U1209/U1125/U28/U1/U2  ( .x(\U1209/U1125/U28/U1/set ), .a(xsel), 
        .b(\U1209/nack[1] ), .c(\U1209/nack[0] ) );
    nand2_2 \U1209/U1125/U28/U1/U3  ( .x(nxa), .a(\U1209/U1125/U28/U1/clr ), 
        .b(\U1209/U1125/U28/U1/set ) );
    aoai211_1 \U1209/U1122/U28/U1/U1  ( .x(\U1209/U1122/U28/U1/clr ), .a(
        \U1209/nack[0] ), .b(\U1209/nack[1] ), .c(ysel), .d(nyla) );
    nand3_1 \U1209/U1122/U28/U1/U2  ( .x(\U1209/U1122/U28/U1/set ), .a(ysel), 
        .b(\U1209/nack[0] ), .c(\U1209/nack[1] ) );
    nand2_2 \U1209/U1122/U28/U1/U3  ( .x(nyla), .a(\U1209/U1122/U28/U1/clr ), 
        .b(\U1209/U1122/U28/U1/set ) );
    oa31_1 \U1209/U916_0_/U25/U1/Uclr  ( .x(\U1209/U916_0_/U25/U1/clr ), .a(
        noa), .b(\x[0] ), .c(\yl[0] ), .d(o[0]) );
    oaoi211_1 \U1209/U916_0_/U25/U1/Uaoi  ( .x(\U1209/U916_0_/U25/U1/ob ), .a(
        \x[0] ), .b(\yl[0] ), .c(noa), .d(\U1209/U916_0_/U25/U1/clr ) );
    inv_2 \U1209/U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U1209/U916_0_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_1_/U25/U1/Uclr  ( .x(\U1209/U916_1_/U25/U1/clr ), .a(
        noa), .b(\x[1] ), .c(\yl[1] ), .d(o[1]) );
    oaoi211_1 \U1209/U916_1_/U25/U1/Uaoi  ( .x(\U1209/U916_1_/U25/U1/ob ), .a(
        \x[1] ), .b(\yl[1] ), .c(noa), .d(\U1209/U916_1_/U25/U1/clr ) );
    inv_2 \U1209/U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U1209/U916_1_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_2_/U25/U1/Uclr  ( .x(\U1209/U916_2_/U25/U1/clr ), .a(
        noa), .b(\x[2] ), .c(\yl[2] ), .d(o[2]) );
    oaoi211_1 \U1209/U916_2_/U25/U1/Uaoi  ( .x(\U1209/U916_2_/U25/U1/ob ), .a(
        \x[2] ), .b(\yl[2] ), .c(noa), .d(\U1209/U916_2_/U25/U1/clr ) );
    inv_2 \U1209/U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U1209/U916_2_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_3_/U25/U1/Uclr  ( .x(\U1209/U916_3_/U25/U1/clr ), .a(
        noa), .b(\x[3] ), .c(\yl[3] ), .d(o[3]) );
    oaoi211_1 \U1209/U916_3_/U25/U1/Uaoi  ( .x(\U1209/U916_3_/U25/U1/ob ), .a(
        \x[3] ), .b(\yl[3] ), .c(noa), .d(\U1209/U916_3_/U25/U1/clr ) );
    inv_2 \U1209/U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U1209/U916_3_/U25/U1/ob )
         );
    nor2_1 \U1213/U1128/U5  ( .x(\U1213/nack[0] ), .a(\y[3] ), .b(\y[2] ) );
    nor3_1 \U1213/U1127/U7  ( .x(\U1213/nack[1] ), .a(\y[1] ), .b(\U1213/net4 
        ), .c(\y[0] ) );
    inv_1 \U1213/U907/U3  ( .x(\U1213/net4 ), .a(nbReset) );
    aoai211_1 \U1213/U1125/U28/U1/U1  ( .x(\U1213/U1125/U28/U1/clr ), .a(
        \U1213/nack[1] ), .b(\U1213/nack[0] ), .c(bsel), .d(nba) );
    nand3_1 \U1213/U1125/U28/U1/U2  ( .x(\U1213/U1125/U28/U1/set ), .a(bsel), 
        .b(\U1213/nack[1] ), .c(\U1213/nack[0] ) );
    nand2_2 \U1213/U1125/U28/U1/U3  ( .x(nba), .a(\U1213/U1125/U28/U1/clr ), 
        .b(\U1213/U1125/U28/U1/set ) );
    aoai211_1 \U1213/U1122/U28/U1/U1  ( .x(\U1213/U1122/U28/U1/clr ), .a(
        \U1213/nack[0] ), .b(\U1213/nack[1] ), .c(dsel), .d(nda) );
    nand3_1 \U1213/U1122/U28/U1/U2  ( .x(\U1213/U1122/U28/U1/set ), .a(dsel), 
        .b(\U1213/nack[0] ), .c(\U1213/nack[1] ) );
    nand2_2 \U1213/U1122/U28/U1/U3  ( .x(nda), .a(\U1213/U1122/U28/U1/clr ), 
        .b(\U1213/U1122/U28/U1/set ) );
    oa31_1 \U1213/U916_0_/U25/U1/Uclr  ( .x(\U1213/U916_0_/U25/U1/clr ), .a(
        nya), .b(\b[0] ), .c(\d[0] ), .d(\y[0] ) );
    oaoi211_1 \U1213/U916_0_/U25/U1/Uaoi  ( .x(\U1213/U916_0_/U25/U1/ob ), .a(
        \b[0] ), .b(\d[0] ), .c(nya), .d(\U1213/U916_0_/U25/U1/clr ) );
    inv_2 \U1213/U916_0_/U25/U1/Ui  ( .x(\y[0] ), .a(\U1213/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_1_/U25/U1/Uclr  ( .x(\U1213/U916_1_/U25/U1/clr ), .a(
        nya), .b(\b[1] ), .c(\d[1] ), .d(\y[1] ) );
    oaoi211_1 \U1213/U916_1_/U25/U1/Uaoi  ( .x(\U1213/U916_1_/U25/U1/ob ), .a(
        \b[1] ), .b(\d[1] ), .c(nya), .d(\U1213/U916_1_/U25/U1/clr ) );
    inv_2 \U1213/U916_1_/U25/U1/Ui  ( .x(\y[1] ), .a(\U1213/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_2_/U25/U1/Uclr  ( .x(\U1213/U916_2_/U25/U1/clr ), .a(
        nya), .b(\b[2] ), .c(\d[2] ), .d(\y[2] ) );
    oaoi211_1 \U1213/U916_2_/U25/U1/Uaoi  ( .x(\U1213/U916_2_/U25/U1/ob ), .a(
        \b[2] ), .b(\d[2] ), .c(nya), .d(\U1213/U916_2_/U25/U1/clr ) );
    inv_2 \U1213/U916_2_/U25/U1/Ui  ( .x(\y[2] ), .a(\U1213/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_3_/U25/U1/Uclr  ( .x(\U1213/U916_3_/U25/U1/clr ), .a(
        nya), .b(\b[3] ), .c(\d[3] ), .d(\y[3] ) );
    oaoi211_1 \U1213/U916_3_/U25/U1/Uaoi  ( .x(\U1213/U916_3_/U25/U1/ob ), .a(
        \b[3] ), .b(\d[3] ), .c(nya), .d(\U1213/U916_3_/U25/U1/clr ) );
    inv_2 \U1213/U916_3_/U25/U1/Ui  ( .x(\y[3] ), .a(\U1213/U916_3_/U25/U1/ob 
        ) );
    and3_2 \U1210/U1138/U9  ( .x(\d[3] ), .a(\cdh[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1137/U9  ( .x(\d[2] ), .a(\cdl[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1139/U9  ( .x(\d[1] ), .a(\cdh[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1210/U1136/U9  ( .x(\d[0] ), .a(\cdl[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1162/U1138/U9  ( .x(\a[3] ), .a(ih[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1137/U9  ( .x(\a[2] ), .a(il[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1139/U9  ( .x(\a[1] ), .a(ih[6]), .b(naa), .c(il[7]) );
    and3_2 \U1162/U1136/U9  ( .x(\a[0] ), .a(il[6]), .b(naa), .c(il[7]) );
    and3_2 \U1211/U1138/U9  ( .x(\b[3] ), .a(ih[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1137/U9  ( .x(\b[2] ), .a(il[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1139/U9  ( .x(\b[1] ), .a(ih[4]), .b(nba), .c(il[5]) );
    and3_2 \U1211/U1136/U9  ( .x(\b[0] ), .a(il[4]), .b(nba), .c(il[5]) );
    and3_2 \U1163/U1138/U9  ( .x(\c[3] ), .a(\cdh[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1137/U9  ( .x(\c[2] ), .a(\cdl[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1139/U9  ( .x(\c[1] ), .a(\cdh[2] ), .b(nca), .c(\cdl[3] )
         );
    and3_2 \U1163/U1136/U9  ( .x(\c[0] ), .a(\cdl[2] ), .b(nca), .c(\cdl[3] )
         );
    and2_1 \U1296/U1385/U8  ( .x(cg), .a(nbReset), .b(\U1296/ng ) );
    aoi222_1 \U1296/U1384/U30/U1  ( .x(\U1296/ng ), .a(nca), .b(net195), .c(
        nca), .d(\U1296/U1384/Z ), .e(net195), .f(\U1296/U1384/Z ) );
    inv_1 \U1296/U1384/U30/Uinv  ( .x(\U1296/U1384/Z ), .a(\U1296/ng ) );
    oa31_1 \U1296/U1386/U25/U1/Uclr  ( .x(\U1296/U1386/U25/U1/clr ), .a(
        \twobitack[2] ), .b(cg), .c(nca), .d(net195) );
    oaoi211_1 \U1296/U1386/U25/U1/Uaoi  ( .x(\U1296/U1386/U25/U1/ob ), .a(cg), 
        .b(nca), .c(\twobitack[2] ), .d(\U1296/U1386/U25/U1/clr ) );
    inv_2 \U1296/U1386/U25/U1/Ui  ( .x(net195), .a(\U1296/U1386/U25/U1/ob ) );
    and2_1 \U1298/U1385/U8  ( .x(dg), .a(nbReset), .b(\U1298/ng ) );
    aoi222_1 \U1298/U1384/U30/U1  ( .x(\U1298/ng ), .a(nda), .b(net193), .c(
        nda), .d(\U1298/U1384/Z ), .e(net193), .f(\U1298/U1384/Z ) );
    inv_1 \U1298/U1384/U30/Uinv  ( .x(\U1298/U1384/Z ), .a(\U1298/ng ) );
    oa31_1 \U1298/U1386/U25/U1/Uclr  ( .x(\U1298/U1386/U25/U1/clr ), .a(
        \twobitack[0] ), .b(dg), .c(nda), .d(net193) );
    oaoi211_1 \U1298/U1386/U25/U1/Uaoi  ( .x(\U1298/U1386/U25/U1/ob ), .a(dg), 
        .b(nda), .c(\twobitack[0] ), .d(\U1298/U1386/U25/U1/clr ) );
    inv_2 \U1298/U1386/U25/U1/Ui  ( .x(net193), .a(\U1298/U1386/U25/U1/ob ) );
    and2_1 \U1306/U1385/U8  ( .x(bg), .a(nbReset), .b(\U1306/ng ) );
    aoi222_1 \U1306/U1384/U30/U1  ( .x(\U1306/ng ), .a(nba), .b(\twobitack[1] 
        ), .c(nba), .d(\U1306/U1384/Z ), .e(\twobitack[1] ), .f(
        \U1306/U1384/Z ) );
    inv_1 \U1306/U1384/U30/Uinv  ( .x(\U1306/U1384/Z ), .a(\U1306/ng ) );
    oa31_1 \U1306/U1386/U25/U1/Uclr  ( .x(\U1306/U1386/U25/U1/clr ), .a(net199
        ), .b(bg), .c(nba), .d(\twobitack[1] ) );
    oaoi211_1 \U1306/U1386/U25/U1/Uaoi  ( .x(\U1306/U1386/U25/U1/ob ), .a(bg), 
        .b(nba), .c(net199), .d(\U1306/U1386/U25/U1/clr ) );
    inv_2 \U1306/U1386/U25/U1/Ui  ( .x(\twobitack[1] ), .a(
        \U1306/U1386/U25/U1/ob ) );
    and2_1 \U1295/U1385/U8  ( .x(ag), .a(nbReset), .b(\U1295/ng ) );
    aoi222_1 \U1295/U1384/U30/U1  ( .x(\U1295/ng ), .a(naa), .b(\twobitack[3] 
        ), .c(naa), .d(\U1295/U1384/Z ), .e(\twobitack[3] ), .f(
        \U1295/U1384/Z ) );
    inv_1 \U1295/U1384/U30/Uinv  ( .x(\U1295/U1384/Z ), .a(\U1295/ng ) );
    oa31_1 \U1295/U1386/U25/U1/Uclr  ( .x(\U1295/U1386/U25/U1/clr ), .a(net194
        ), .b(ag), .c(naa), .d(\twobitack[3] ) );
    oaoi211_1 \U1295/U1386/U25/U1/Uaoi  ( .x(\U1295/U1386/U25/U1/ob ), .a(ag), 
        .b(naa), .c(net194), .d(\U1295/U1386/U25/U1/clr ) );
    inv_2 \U1295/U1386/U25/U1/Ui  ( .x(\twobitack[3] ), .a(
        \U1295/U1386/U25/U1/ob ) );
    nand2_1 \U1297/U1131/U5  ( .x(\U1297/s ), .a(\U1297/r ), .b(\U1297/nback )
         );
    nand2_1 \U1297/U1103/U5  ( .x(\U1297/r ), .a(\U1297/naack ), .b(\U1297/s )
         );
    inv_1 \U1297/U1111/U3  ( .x(\U1297/reset ), .a(nbReset) );
    inv_1 \U1297/U1112/U3  ( .x(\U1297/naack ), .a(naa) );
    nor2_1 \U1297/U1130/U5  ( .x(\U1297/nback ), .a(nca), .b(\U1297/reset ) );
    aoai211_1 \U1297/U1128/U28/U1/U1  ( .x(\U1297/U1128/U28/U1/clr ), .a(
        \U1297/r ), .b(\U1297/naack ), .c(cg), .d(csel) );
    nand3_1 \U1297/U1128/U28/U1/U2  ( .x(\U1297/U1128/U28/U1/set ), .a(cg), 
        .b(\U1297/r ), .c(\U1297/naack ) );
    nand2_2 \U1297/U1128/U28/U1/U3  ( .x(csel), .a(\U1297/U1128/U28/U1/clr ), 
        .b(\U1297/U1128/U28/U1/set ) );
    aoai211_1 \U1297/U1127/U28/U1/U1  ( .x(\U1297/U1127/U28/U1/clr ), .a(
        \U1297/s ), .b(\U1297/nback ), .c(ag), .d(asel) );
    nand3_1 \U1297/U1127/U28/U1/U2  ( .x(\U1297/U1127/U28/U1/set ), .a(ag), 
        .b(\U1297/s ), .c(\U1297/nback ) );
    nand2_2 \U1297/U1127/U28/U1/U3  ( .x(asel), .a(\U1297/U1127/U28/U1/clr ), 
        .b(\U1297/U1127/U28/U1/set ) );
    nand2_1 \U1300/U1131/U5  ( .x(\U1300/s ), .a(\U1300/r ), .b(\U1300/nback )
         );
    nand2_1 \U1300/U1103/U5  ( .x(\U1300/r ), .a(\U1300/naack ), .b(\U1300/s )
         );
    inv_1 \U1300/U1111/U3  ( .x(\U1300/reset ), .a(nbReset) );
    inv_1 \U1300/U1112/U3  ( .x(\U1300/naack ), .a(nba) );
    nor2_1 \U1300/U1130/U5  ( .x(\U1300/nback ), .a(nda), .b(\U1300/reset ) );
    aoai211_1 \U1300/U1128/U28/U1/U1  ( .x(\U1300/U1128/U28/U1/clr ), .a(
        \U1300/r ), .b(\U1300/naack ), .c(dg), .d(dsel) );
    nand3_1 \U1300/U1128/U28/U1/U2  ( .x(\U1300/U1128/U28/U1/set ), .a(dg), 
        .b(\U1300/r ), .c(\U1300/naack ) );
    nand2_2 \U1300/U1128/U28/U1/U3  ( .x(dsel), .a(\U1300/U1128/U28/U1/clr ), 
        .b(\U1300/U1128/U28/U1/set ) );
    aoai211_1 \U1300/U1127/U28/U1/U1  ( .x(\U1300/U1127/U28/U1/clr ), .a(
        \U1300/s ), .b(\U1300/nback ), .c(bg), .d(bsel) );
    nand3_1 \U1300/U1127/U28/U1/U2  ( .x(\U1300/U1127/U28/U1/set ), .a(bg), 
        .b(\U1300/s ), .c(\U1300/nback ) );
    nand2_2 \U1300/U1127/U28/U1/U3  ( .x(bsel), .a(\U1300/U1127/U28/U1/clr ), 
        .b(\U1300/U1127/U28/U1/set ) );
    aoai211_1 \U1289/U1150/U28/U1/U1  ( .x(\U1289/U1150/U28/U1/clr ), .a(il[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[2] ) );
    nand3_1 \U1289/U1150/U28/U1/U2  ( .x(\U1289/U1150/U28/U1/set ), .a(net195), 
        .b(il[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1150/U28/U1/U3  ( .x(\cdl[2] ), .a(
        \U1289/U1150/U28/U1/clr ), .b(\U1289/U1150/U28/U1/set ) );
    aoai211_1 \U1289/U1152/U28/U1/U1  ( .x(\U1289/U1152/U28/U1/clr ), .a(il[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[3] ) );
    nand3_1 \U1289/U1152/U28/U1/U2  ( .x(\U1289/U1152/U28/U1/set ), .a(net195), 
        .b(il[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1152/U28/U1/U3  ( .x(\cdl[3] ), .a(
        \U1289/U1152/U28/U1/clr ), .b(\U1289/U1152/U28/U1/set ) );
    aoai211_1 \U1289/U1149/U28/U1/U1  ( .x(\U1289/U1149/U28/U1/clr ), .a(ih[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[2] ) );
    nand3_1 \U1289/U1149/U28/U1/U2  ( .x(\U1289/U1149/U28/U1/set ), .a(net195), 
        .b(ih[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1149/U28/U1/U3  ( .x(\cdh[2] ), .a(
        \U1289/U1149/U28/U1/clr ), .b(\U1289/U1149/U28/U1/set ) );
    aoai211_1 \U1289/U1151/U28/U1/U1  ( .x(\U1289/U1151/U28/U1/clr ), .a(ih[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[3] ) );
    nand3_1 \U1289/U1151/U28/U1/U2  ( .x(\U1289/U1151/U28/U1/set ), .a(net195), 
        .b(ih[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1151/U28/U1/U3  ( .x(\cdh[3] ), .a(
        \U1289/U1151/U28/U1/clr ), .b(\U1289/U1151/U28/U1/set ) );
    inv_1 \U1289/U1148/U1147/U3  ( .x(\U1289/U1148/net189 ), .a(
        \U1289/bnreset ) );
    nor2_1 \U1289/U1148/U582/U5  ( .x(\U1289/U1148/net192 ), .a(\cdl[3] ), .b(
        \cdh[3] ) );
    nor2_1 \U1289/U1148/U580/U5  ( .x(\U1289/U1148/net191 ), .a(\cdl[2] ), .b(
        \cdh[2] ) );
    nor2_2 \U1289/U1148/U1146/U6  ( .x(\twobitack[2] ), .a(
        \U1289/U1148/net190 ), .b(\U1289/U1148/net189 ) );
    aoi222_1 \U1289/U1148/U1141/U30/U1  ( .x(\U1289/U1148/net190 ), .a(
        \U1289/U1148/net191 ), .b(\U1289/U1148/net192 ), .c(
        \U1289/U1148/net191 ), .d(\U1289/U1148/U1141/Z ), .e(
        \U1289/U1148/net192 ), .f(\U1289/U1148/U1141/Z ) );
    inv_1 \U1289/U1148/U1141/U30/Uinv  ( .x(\U1289/U1148/U1141/Z ), .a(
        \U1289/U1148/net190 ) );
    aoai211_1 \U1271/U1150/U28/U1/U1  ( .x(\U1271/U1150/U28/U1/clr ), .a(il[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[0] ) );
    nand3_1 \U1271/U1150/U28/U1/U2  ( .x(\U1271/U1150/U28/U1/set ), .a(net193), 
        .b(il[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1150/U28/U1/U3  ( .x(\cdl[0] ), .a(
        \U1271/U1150/U28/U1/clr ), .b(\U1271/U1150/U28/U1/set ) );
    aoai211_1 \U1271/U1152/U28/U1/U1  ( .x(\U1271/U1152/U28/U1/clr ), .a(il[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[1] ) );
    nand3_1 \U1271/U1152/U28/U1/U2  ( .x(\U1271/U1152/U28/U1/set ), .a(net193), 
        .b(il[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1152/U28/U1/U3  ( .x(\cdl[1] ), .a(
        \U1271/U1152/U28/U1/clr ), .b(\U1271/U1152/U28/U1/set ) );
    aoai211_1 \U1271/U1149/U28/U1/U1  ( .x(\U1271/U1149/U28/U1/clr ), .a(ih[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[0] ) );
    nand3_1 \U1271/U1149/U28/U1/U2  ( .x(\U1271/U1149/U28/U1/set ), .a(net193), 
        .b(ih[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1149/U28/U1/U3  ( .x(\cdh[0] ), .a(
        \U1271/U1149/U28/U1/clr ), .b(\U1271/U1149/U28/U1/set ) );
    aoai211_1 \U1271/U1151/U28/U1/U1  ( .x(\U1271/U1151/U28/U1/clr ), .a(ih[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[1] ) );
    nand3_1 \U1271/U1151/U28/U1/U2  ( .x(\U1271/U1151/U28/U1/set ), .a(net193), 
        .b(ih[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1151/U28/U1/U3  ( .x(\cdh[1] ), .a(
        \U1271/U1151/U28/U1/clr ), .b(\U1271/U1151/U28/U1/set ) );
    inv_1 \U1271/U1148/U1147/U3  ( .x(\U1271/U1148/net189 ), .a(
        \U1271/bnreset ) );
    nor2_1 \U1271/U1148/U582/U5  ( .x(\U1271/U1148/net192 ), .a(\cdl[1] ), .b(
        \cdh[1] ) );
    nor2_1 \U1271/U1148/U580/U5  ( .x(\U1271/U1148/net191 ), .a(\cdl[0] ), .b(
        \cdh[0] ) );
    nor2_2 \U1271/U1148/U1146/U6  ( .x(\twobitack[0] ), .a(
        \U1271/U1148/net190 ), .b(\U1271/U1148/net189 ) );
    aoi222_1 \U1271/U1148/U1141/U30/U1  ( .x(\U1271/U1148/net190 ), .a(
        \U1271/U1148/net191 ), .b(\U1271/U1148/net192 ), .c(
        \U1271/U1148/net191 ), .d(\U1271/U1148/U1141/Z ), .e(
        \U1271/U1148/net192 ), .f(\U1271/U1148/U1141/Z ) );
    inv_1 \U1271/U1148/U1141/U30/Uinv  ( .x(\U1271/U1148/U1141/Z ), .a(
        \U1271/U1148/net190 ) );
    nand2_1 \U1225/U1128/U5  ( .x(\U1225/s ), .a(\U1225/r ), .b(\U1225/nback )
         );
    nand2_1 \U1225/U1103/U5  ( .x(\U1225/r ), .a(\U1225/naack ), .b(\U1225/s )
         );
    inv_1 \U1225/U1111/U3  ( .x(\U1225/reset ), .a(nbReset) );
    inv_1 \U1225/U1112/U3  ( .x(\U1225/naack ), .a(nxa) );
    nor2_1 \U1225/U1127/U5  ( .x(\U1225/nback ), .a(nyla), .b(\U1225/reset )
         );
    and2_2 \U1225/U1129/U8  ( .x(xsel), .a(\U1225/nback ), .b(\U1225/s ) );
    and2_2 \U1225/U1124/U8  ( .x(ysel), .a(\U1225/r ), .b(\U1225/naack ) );
    and3_4 \U1308/U20/U9  ( .x(nya), .a(\U1308/nack[1] ), .b(\U1308/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U1308/U18/U5  ( .x(\U1308/nack[0] ), .a(\yl[3] ), .b(\yl[0] ) );
    nor2_1 \U1308/U19/U5  ( .x(\U1308/nack[1] ), .a(\yl[1] ), .b(\yl[2] ) );
    ao222_2 \U1308/U15_0_/U19/U1/U1  ( .x(\yl[0] ), .a(\y[0] ), .b(nyla), .c(
        \y[0] ), .d(\yl[0] ), .e(nyla), .f(\yl[0] ) );
    ao222_2 \U1308/U15_1_/U19/U1/U1  ( .x(\yl[1] ), .a(\y[1] ), .b(nyla), .c(
        \y[1] ), .d(\yl[1] ), .e(nyla), .f(\yl[1] ) );
    ao222_2 \U1308/U15_2_/U19/U1/U1  ( .x(\yl[2] ), .a(\y[2] ), .b(nyla), .c(
        \y[2] ), .d(\yl[2] ), .e(nyla), .f(\yl[2] ) );
    ao222_2 \U1308/U15_3_/U19/U1/U1  ( .x(\yl[3] ), .a(\y[3] ), .b(nyla), .c(
        \y[3] ), .d(\yl[3] ), .e(nyla), .f(\yl[3] ) );
    buf_3 U1 ( .x(\U1271/bnreset ), .a(nbReset) );
    buf_3 U2 ( .x(\U1289/bnreset ), .a(nbReset) );
endmodule


module chain_dr8bit_completion_40 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_41 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_42 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_43 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr32bit_completion_9 ( o, i );
input  [63:0] i;
output o;
    wire nx, \cd[3] , \cd[2] , ny, \cd[0] , \cd[1] , \U16/Z , \U6/Z , \U15/Z ;
    chain_dr8bit_completion_40 U11 ( .o(\cd[3] ), .i({i[63], i[62], i[61], 
        i[60], i[59], i[58], i[57], i[56], i[31], i[30], i[29], i[28], i[27], 
        i[26], i[25], i[24]}) );
    chain_dr8bit_completion_43 U14 ( .o(\cd[2] ), .i({i[55], i[54], i[53], 
        i[52], i[51], i[50], i[49], i[48], i[23], i[22], i[21], i[20], i[19], 
        i[18], i[17], i[16]}) );
    chain_dr8bit_completion_42 U13 ( .o(\cd[1] ), .i({i[47], i[46], i[45], 
        i[44], i[43], i[42], i[41], i[40], i[15], i[14], i[13], i[12], i[11], 
        i[10], i[9], i[8]}) );
    chain_dr8bit_completion_41 U12 ( .o(\cd[0] ), .i({i[39], i[38], i[37], 
        i[36], i[35], i[34], i[33], i[32], i[7], i[6], i[5], i[4], i[3], i[2], 
        i[1], i[0]}) );
    aoi222_1 \U16/U30/U1  ( .x(ny), .a(\cd[0] ), .b(\cd[1] ), .c(\cd[0] ), .d(
        \U16/Z ), .e(\cd[1] ), .f(\U16/Z ) );
    inv_1 \U16/U30/Uinv  ( .x(\U16/Z ), .a(ny) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(ny), .b(nx), .c(ny), .d(\U6/Z ), .e(nx), 
        .f(\U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U15/U30/U1  ( .x(nx), .a(\cd[3] ), .b(\cd[2] ), .c(\cd[3] ), .d(
        \U15/Z ), .e(\cd[2] ), .f(\U15/Z ) );
    inv_1 \U15/U30/Uinv  ( .x(\U15/Z ), .a(nx) );
endmodule


module chain_selement_ga_70 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_71 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_t_ctrl_1 ( cack, fcdefer, fcslowack, screq, ack, defer, fcack, 
    nReset, scack, slowack );
input  ack, defer, fcack, nReset, scack, slowack;
output cack, fcdefer, fcslowack, screq;
    wire net269, net280, net275, net270, net265, net278, net276, net277, 
        net263, net271, net266, net279, net272, net264, net267, net273, net268, 
        net274, \U49/U28/U1/clr , \U49/U28/U1/set , \U50/U28/U1/clr , 
        \U50/U28/U1/set , \U51/U28/U1/clr , \U51/U28/U1/set , \U57/acb , 
        \U57/U1/Z ;
    chain_selement_ga_71 U55 ( .Aa(net269), .Br(fcdefer), .Ar(net280), .Ba(
        fcack) );
    chain_selement_ga_70 U54 ( .Aa(net275), .Br(fcslowack), .Ar(net270), .Ba(
        fcack) );
    or2_4 \U12/U12  ( .x(net268), .a(net266), .b(net270) );
    or2_4 \U56/U12  ( .x(net274), .a(net275), .b(net269) );
    or2_4 \U14/U12  ( .x(net273), .a(net274), .b(net266) );
    or3_1 \U36/U12  ( .x(cack), .a(net267), .b(net264), .c(net272) );
    nor3_1 \U21/U7  ( .x(net271), .a(net270), .b(net266), .c(net280) );
    and2_1 \U53/U8  ( .x(net263), .a(net271), .b(nReset) );
    and2_1 \U43/U8  ( .x(net277), .a(net265), .b(nReset) );
    nor2_1 \U22/U5  ( .x(net265), .a(net278), .b(net276) );
    ao222_2 \U44/U19/U1/U1  ( .x(net276), .a(net280), .b(net273), .c(net280), 
        .d(net276), .e(net273), .f(net276) );
    ao222_2 \U40/U19/U1/U1  ( .x(net280), .a(net272), .b(net277), .c(net272), 
        .d(net280), .e(net277), .f(net280) );
    ao222_2 \U45/U19/U1/U1  ( .x(net279), .a(net273), .b(net268), .c(net273), 
        .d(net279), .e(net268), .f(net279) );
    ao222_2 \U42/U19/U1/U1  ( .x(net266), .a(net277), .b(net267), .c(net277), 
        .d(net266), .e(net267), .f(net266) );
    ao222_2 \U39/U19/U1/U1  ( .x(net270), .a(net277), .b(net264), .c(net277), 
        .d(net270), .e(net264), .f(net270) );
    aoai211_1 \U49/U28/U1/U1  ( .x(\U49/U28/U1/clr ), .a(ack), .b(nReset), .c(
        net263), .d(net267) );
    nand3_1 \U49/U28/U1/U2  ( .x(\U49/U28/U1/set ), .a(net263), .b(ack), .c(
        nReset) );
    nand2_2 \U49/U28/U1/U3  ( .x(net267), .a(\U49/U28/U1/clr ), .b(
        \U49/U28/U1/set ) );
    aoai211_1 \U50/U28/U1/U1  ( .x(\U50/U28/U1/clr ), .a(slowack), .b(nReset), 
        .c(net263), .d(net264) );
    nand3_1 \U50/U28/U1/U2  ( .x(\U50/U28/U1/set ), .a(net263), .b(slowack), 
        .c(nReset) );
    nand2_2 \U50/U28/U1/U3  ( .x(net264), .a(\U50/U28/U1/clr ), .b(
        \U50/U28/U1/set ) );
    aoai211_1 \U51/U28/U1/U1  ( .x(\U51/U28/U1/clr ), .a(defer), .b(nReset), 
        .c(net263), .d(net272) );
    nand2_2 \U51/U28/U1/U3  ( .x(net272), .a(\U51/U28/U1/clr ), .b(
        \U51/U28/U1/set ) );
    and2_1 \U57/U2/U8  ( .x(screq), .a(net279), .b(\U57/acb ) );
    nor2_1 \U57/U3/U5  ( .x(net278), .a(\U57/acb ), .b(scack) );
    oai21_1 \U57/U1/U30/U1/U1  ( .x(\U57/acb ), .a(\U57/U1/Z ), .b(scack), .c(
        net279) );
    inv_1 \U57/U1/U30/U1/U2  ( .x(\U57/U1/Z ), .a(\U57/acb ) );
    nand3_0 U1 ( .x(\U51/U28/U1/set ), .a(net263), .b(defer), .c(nReset) );
endmodule


module chain_mergepackets_4 ( naa, nba, o, a, b, nReset, noa );
output [4:0] o;
input  [4:0] a;
input  [4:0] b;
input  nReset, noa;
output naa, nba;
    wire \noack[1] , \noack[0] , reset, bsel, as, setb, asel, seta, 
        \U916_0_/U25/U1/clr , \U916_0_/U25/U1/ob , \U916_1_/U25/U1/clr , 
        \U916_1_/U25/U1/ob , \U916_2_/U25/U1/clr , \U916_2_/U25/U1/ob , 
        \U916_3_/U25/U1/clr , \U916_3_/U25/U1/ob ;
    and2_1 \U1155/U8  ( .x(as), .a(seta), .b(asel) );
    nand2_1 \U1145/U5  ( .x(asel), .a(bsel), .b(seta) );
    nand2_1 \U1103/U5  ( .x(bsel), .a(setb), .b(asel) );
    inv_1 \U1135/U3  ( .x(reset), .a(nReset) );
    inv_1 \U1134/U3  ( .x(setb), .a(a[4]) );
    and3_2 \U1154/U9  ( .x(naa), .a(\noack[1] ), .b(\noack[0] ), .c(as) );
    nor3_1 \U1127/U7  ( .x(\noack[0] ), .a(o[1]), .b(reset), .c(o[0]) );
    nor2_1 \U1132/U5  ( .x(\noack[1] ), .a(o[3]), .b(o[2]) );
    oa31_1 \U916_0_/U25/U1/Uclr  ( .x(\U916_0_/U25/U1/clr ), .a(noa), .b(a[0]), 
        .c(b[0]), .d(o[0]) );
    oaoi211_1 \U916_0_/U25/U1/Uaoi  ( .x(\U916_0_/U25/U1/ob ), .a(a[0]), .b(b
        [0]), .c(noa), .d(\U916_0_/U25/U1/clr ) );
    inv_2 \U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U916_0_/U25/U1/ob ) );
    oa31_1 \U916_1_/U25/U1/Uclr  ( .x(\U916_1_/U25/U1/clr ), .a(noa), .b(a[1]), 
        .c(b[1]), .d(o[1]) );
    oaoi211_1 \U916_1_/U25/U1/Uaoi  ( .x(\U916_1_/U25/U1/ob ), .a(a[1]), .b(b
        [1]), .c(noa), .d(\U916_1_/U25/U1/clr ) );
    inv_2 \U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U916_1_/U25/U1/ob ) );
    oa31_1 \U916_2_/U25/U1/Uclr  ( .x(\U916_2_/U25/U1/clr ), .a(noa), .b(a[2]), 
        .c(b[2]), .d(o[2]) );
    oaoi211_1 \U916_2_/U25/U1/Uaoi  ( .x(\U916_2_/U25/U1/ob ), .a(a[2]), .b(b
        [2]), .c(noa), .d(\U916_2_/U25/U1/clr ) );
    inv_2 \U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U916_2_/U25/U1/ob ) );
    oa31_1 \U916_3_/U25/U1/Uclr  ( .x(\U916_3_/U25/U1/clr ), .a(noa), .b(a[3]), 
        .c(b[3]), .d(o[3]) );
    oaoi211_1 \U916_3_/U25/U1/Uaoi  ( .x(\U916_3_/U25/U1/ob ), .a(a[3]), .b(b
        [3]), .c(noa), .d(\U916_3_/U25/U1/clr ) );
    inv_2 \U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U916_3_/U25/U1/ob ) );
    ao222_2 \U1148/U19/U1/U1  ( .x(o[4]), .a(noa), .b(b[4]), .c(noa), .d(o[4]), 
        .e(b[4]), .f(o[4]) );
    aoi21_1 \U1153/U11  ( .x(seta), .a(o[4]), .b(setb), .c(reset) );
    and3_3 U1 ( .x(nba), .a(bsel), .b(\noack[0] ), .c(\noack[1] ) );
endmodule


module target_imem ( addr, ccol, chainresponse, crnw, csize, ctag, lock, 
    nchaincommandack, nrouteack, pred, rack, routetxreq, seq, tag_h, tag_l, wd, 
    cack, cdefer, chaincommand, cndefer, cok, err, nReset, nchainresponseack, 
    rd, route, routetxack );
output [63:0] addr;
output [5:0] ccol;
output [4:0] chainresponse;
output [1:0] crnw;
output [3:0] csize;
output [9:0] ctag;
output [1:0] lock;
output [1:0] pred;
output [1:0] seq;
output [4:0] tag_h;
output [4:0] tag_l;
output [63:0] wd;
input  [4:0] chaincommand;
input  [1:0] err;
input  [63:0] rd;
input  [4:0] route;
input  cack, cdefer, cndefer, cok, nReset, nchainresponseack, routetxack;
output nchaincommandack, nrouteack, rack, routetxreq;
    wire n9, n10, n11, n12, \net242[0] , \net242[1] , \net242[2] , \net242[3] , 
        \net242[4] , \net242[5] , \net242[6] , \net242[7] , \net242[8] , 
        \net242[9] , \net242[10] , \net243[0] , \net243[1] , \net243[2] , 
        \net243[3] , \net243[4] , \net243[5] , \net243[6] , \net243[7] , 
        \net243[8] , \net243[9] , \net243[10] , \net244[0] , \net244[1] , 
        \net244[2] , \net244[3] , \net244[4] , \net244[5] , \net244[6] , 
        \net244[7] , \net244[8] , \net244[9] , \net244[10] , \chainff_l[7] , 
        \chainff_l[6] , \chainff_l[5] , \chainff_l[4] , \chainff_l[3] , 
        \chainff_l[2] , \chainff_l[1] , \chainff_l[0] , \chdrack[0] , 
        \chdrack[1] , \obl[7] , \obl[6] , \obl[5] , \obl[4] , \obl[3] , 
        \obl[2] , \obl[1] , \obl[0] , \tcbh[7] , \tcbh[6] , \tcbh[5] , 
        \tcbh[4] , \tcbh[3] , \tcbh[2] , \tcbh[1] , \tcbh[0] , \tcbl[7] , 
        \tcbl[6] , \tcbl[5] , \tcbl[4] , \tcbl[3] , \tcbl[2] , \tcbl[1] , 
        \tcbl[0] , \tresponse[4] , \tresponse[3] , \tresponse[2] , 
        \tresponse[1] , \tresponse[0] , \nchdr_ack[10] , \nchdr_ack[9] , 
        \nchdr_ack[8] , \nchdr_ack[7] , \nchdr_ack[6] , \nchdr_ack[5] , 
        \nchdr_ack[4] , \nchdr_ack[3] , \nchdr_ack[2] , \nchdr_ack[1] , 
        \nchdr_ack[0] , \chainff_h[7] , \chainff_h[6] , \chainff_h[5] , 
        \chainff_h[4] , \chainff_h[3] , \chainff_h[2] , \chainff_h[1] , 
        \chainff_h[0] , \rhdr_l[15] , \rhdr_l[14] , \rhdr_l[13] , \rhdr_l[7] , 
        \rhdr_l[6] , \rhdr_l[5] , \obh[7] , \obh[6] , \obh[5] , \obh[4] , 
        \obh[3] , \obh[2] , \obh[1] , \obh[0] , \rhdr_h[15] , \rhdr_h[14] , 
        \rhdr_h[13] , \rhdr_h[7] , \rhdr_h[6] , \rhdr_h[5] , net265, nbreset, 
        net248, rhdrack, read_ctrlack, chainff_ack, read_req, read_cd, teop, 
        fcack, tcba, net145, screq, fcslowack, fcdefer, read_ack, 
        ntresponseack, net200, noba, pullcd, net168, net188, net201, net194, 
        net178, net189, net191, net284, hdrcd, chdrctrlack, \U1770/U21/nr , 
        \U1770/U21/nd , \U1770/U21/n2 , \U1761/U28/Z , \U1761/U32/Z , 
        \U1761/U29/Z , \U1761/U33/Z , \U1761/U30/Z , \U1761/U31/Z , \U1632/Z , 
        \U1676/Z , \U1761/y[0] , \U1761/y[1] , \U1761/x[1] , \U1761/x[3] , 
        \U1761/x[2] , \U1761/x[0] , \U1574_0_/net231 , \U1574_1_/net231 , 
        \U1574_2_/net231 , \U1574_3_/net231 , \U1574_4_/net231 , 
        \U1574_5_/net231 , \U1574_6_/net231 , \U1574_7_/net231 , 
        \U1574_8_/net231 , \U1574_9_/net231 , \U1574_10_/net231 , n5, n6, n7, 
        n8;
    chain_sendword_1 U1765 ( .ctrlack(read_ctrlack), .oh({\chainff_h[7] , 
        \chainff_h[6] , \chainff_h[5] , \chainff_h[4] , \chainff_h[3] , 
        \chainff_h[2] , \chainff_h[1] , \chainff_h[0] }), .ol({\chainff_l[7] , 
        \chainff_l[6] , \chainff_l[5] , \chainff_l[4] , \chainff_l[3] , 
        \chainff_l[2] , \chainff_l[1] , \chainff_l[0] }), .chainackff(
        chainff_ack), .ctrlreq(read_req), .ih(rd[63:32]), .il(rd[31:0]) );
    chain_dr32bit_completion_9 rd_cd ( .o(read_cd), .i(rd) );
    chain_trhdr_1 xmitHdr ( .chainff_ack(chainff_ack), .chainh({\tcbh[7] , 
        \tcbh[6] , \tcbh[5] , \tcbh[4] , \tcbh[3] , \tcbh[2] , \tcbh[1] , 
        \tcbh[0] }), .chainl({\tcbl[7] , \tcbl[6] , \tcbl[5] , \tcbl[4] , 
        \tcbl[3] , \tcbl[2] , \tcbl[1] , \tcbl[0] }), .eop(teop), .hdrack(
        rhdrack), .normal_ack(rack), .notify_ack(fcack), .read_req(read_req), 
        .routereq(routetxreq), .chain_ff_h({\chainff_h[7] , \chainff_h[6] , 
        \chainff_h[5] , \chainff_h[4] , \chainff_h[3] , \chainff_h[2] , 
        \chainff_h[1] , \chainff_h[0] }), .chainack(tcba), .chainff_l({
        \chainff_l[7] , \chainff_l[6] , \chainff_l[5] , \chainff_l[4] , 
        \chainff_l[3] , \chainff_l[2] , \chainff_l[1] , \chainff_l[0] }), 
        .eopack(net145), .err(err), .nReset(n5), .normal_response(screq), 
        .notify_accept(fcslowack), .notify_defer(fcdefer), .rcol_h({
        \rhdr_h[15] , \rhdr_h[14] , \rhdr_h[13] }), .rcol_l({\rhdr_l[15] , 
        \rhdr_l[14] , \rhdr_l[13] }), .read_ack(read_ack), .rnw_h(\rhdr_h[7] ), 
        .rnw_l(\rhdr_l[7] ), .routeack(routetxack), .rsize_h({\rhdr_h[6] , 
        \rhdr_h[5] }), .rsize_l({\rhdr_l[6] , \rhdr_l[5] }), .rtag_h(tag_h), 
        .rtag_l(tag_l) );
    chain_dr2fr_byte_4 dr2fr ( .eop_ack(net145), .ia(tcba), .o({\tresponse[4] , 
        \tresponse[3] , \tresponse[2] , \tresponse[1] , \tresponse[0] }), 
        .eop(teop), .ih({\tcbh[7] , \tcbh[6] , \tcbh[5] , \tcbh[4] , \tcbh[3] , 
        \tcbh[2] , \tcbh[1] , \tcbh[0] }), .il({\tcbl[7] , \tcbl[6] , 
        \tcbl[5] , \tcbl[4] , \tcbl[3] , \tcbl[2] , \tcbl[1] , \tcbl[0] }), 
        .nReset(nbreset), .noa(ntresponseack) );
    chain_mergepackets_4 merger ( .naa(nrouteack), .nba(ntresponseack), .o(
        chainresponse), .a(route), .b({\tresponse[4] , \tresponse[3] , 
        \tresponse[2] , \tresponse[1] , \tresponse[0] }), .nReset(nbreset), 
        .noa(nchainresponseack) );
    chain_tchdr_1 header ( .addr_req(net200), .col_h(ccol[5:3]), .col_l(ccol
        [2:0]), .itag_h(ctag[9:5]), .itag_l(ctag[4:0]), .lock(lock), .ncback(
        noba), .pred(pred), .pullcd(pullcd), .reset(net168), .rnw_h(n9), 
        .rnw_l(n10), .seq(seq), .size_h(csize[3:2]), .size_l({n11, n12}), 
        .write_req(net188), .chwh({\obh[7] , \obh[6] , \obh[5] , \obh[4] , 
        \obh[3] , \obh[2] , \obh[1] , \obh[0] }), .chwl({\obl[7] , \obl[6] , 
        \obl[5] , \obl[4] , \obl[3] , \obl[2] , \obl[1] , \obl[0] }), 
        .addr_ack(net201), .addr_pull(net194), .nReset(n5), .nack(net178), 
        .write_ack(net189), .write_pull(net191) );
    chain_irdemux_32new_3 wd_hld ( .ctrlack(net189), .oh(wd[63:32]), .ol(wd
        [31:0]), .pullreq(net191), .pull_h({\obh[7] , \obh[6] , \obh[5] , 
        \obh[4] , \obh[3] , \obh[2] , \obh[1] , \obh[0] }), .pull_l({\obl[7] , 
        \obl[6] , \obl[5] , \obl[4] , \obl[3] , \obl[2] , \obl[1] , \obl[0] }), 
        .pullcd(pullcd), .reset(net168), .ctrlreq(net188) );
    chain_irdemux_32new_2 adr_hld ( .ctrlack(net201), .oh(addr[63:32]), .ol(
        addr[31:0]), .pullreq(net194), .pull_h({\obh[7] , \obh[6] , \obh[5] , 
        \obh[4] , \obh[3] , \obh[2] , \obh[1] , \obh[0] }), .pull_l({\obl[7] , 
        \obl[6] , \obl[5] , \obl[4] , \obl[3] , \obl[2] , \obl[1] , \obl[0] }), 
        .pullcd(pullcd), .reset(net168), .ctrlreq(net200) );
    chain_fr2dr_byte_1 chain_decoder ( .nia(nchaincommandack), .oh({\obh[7] , 
        \obh[6] , \obh[5] , \obh[4] , \obh[3] , \obh[2] , \obh[1] , \obh[0] }), 
        .ol({\obl[7] , \obl[6] , \obl[5] , \obl[4] , \obl[3] , \obl[2] , 
        \obl[1] , \obl[0] }), .i(chaincommand), .nReset(nbreset), .noa(noba)
         );
    chain_t_ctrl_1 cmd_ctrl ( .cack(net284), .fcdefer(fcdefer), .fcslowack(
        fcslowack), .screq(screq), .ack(cok), .defer(cdefer), .fcack(fcack), 
        .nReset(n5), .scack(rack), .slowack(cndefer) );
    inv_1 \I4/U3  ( .x(net265), .a(nbreset) );
    ao222_1 \U1761/U37/U18/U1/U1  ( .x(\chdrack[0] ), .a(\U1761/y[0] ), .b(
        \U1761/y[1] ), .c(\U1761/y[0] ), .d(\chdrack[0] ), .e(\U1761/y[1] ), 
        .f(\chdrack[0] ) );
    ao222_1 \U1762/U18/U1/U1  ( .x(chdrctrlack), .a(hdrcd), .b(net284), .c(
        hdrcd), .d(chdrctrlack), .e(net284), .f(chdrctrlack) );
    ao222_1 \U1769/U18/U1/U1  ( .x(read_ack), .a(read_ctrlack), .b(read_cd), 
        .c(read_ctrlack), .d(read_ack), .e(read_cd), .f(read_ack) );
    aoi222_1 \U1761/U28/U30/U1  ( .x(\U1761/x[3] ), .a(\nchdr_ack[7] ), .b(
        \nchdr_ack[6] ), .c(\nchdr_ack[7] ), .d(\U1761/U28/Z ), .e(
        \nchdr_ack[6] ), .f(\U1761/U28/Z ) );
    inv_1 \U1761/U28/U30/Uinv  ( .x(\U1761/U28/Z ), .a(\U1761/x[3] ) );
    aoi222_1 \U1761/U32/U30/U1  ( .x(\U1761/x[0] ), .a(\nchdr_ack[1] ), .b(
        \nchdr_ack[0] ), .c(\nchdr_ack[1] ), .d(\U1761/U32/Z ), .e(
        \nchdr_ack[0] ), .f(\U1761/U32/Z ) );
    inv_1 \U1761/U32/U30/Uinv  ( .x(\U1761/U32/Z ), .a(\U1761/x[0] ) );
    aoi222_1 \U1761/U29/U30/U1  ( .x(\U1761/x[2] ), .a(\nchdr_ack[5] ), .b(
        \nchdr_ack[4] ), .c(\nchdr_ack[5] ), .d(\U1761/U29/Z ), .e(
        \nchdr_ack[4] ), .f(\U1761/U29/Z ) );
    inv_1 \U1761/U29/U30/Uinv  ( .x(\U1761/U29/Z ), .a(\U1761/x[2] ) );
    aoi222_1 \U1761/U33/U30/U1  ( .x(\U1761/y[0] ), .a(\U1761/x[1] ), .b(
        \U1761/x[0] ), .c(\U1761/x[1] ), .d(\U1761/U33/Z ), .e(\U1761/x[0] ), 
        .f(\U1761/U33/Z ) );
    inv_1 \U1761/U33/U30/Uinv  ( .x(\U1761/U33/Z ), .a(\U1761/y[0] ) );
    aoi222_1 \U1761/U30/U30/U1  ( .x(\U1761/y[1] ), .a(\U1761/x[3] ), .b(
        \U1761/x[2] ), .c(\U1761/x[3] ), .d(\U1761/U30/Z ), .e(\U1761/x[2] ), 
        .f(\U1761/U30/Z ) );
    inv_1 \U1761/U30/U30/Uinv  ( .x(\U1761/U30/Z ), .a(\U1761/y[1] ) );
    aoi222_1 \U1761/U31/U30/U1  ( .x(\U1761/x[1] ), .a(\nchdr_ack[3] ), .b(
        \nchdr_ack[2] ), .c(\nchdr_ack[3] ), .d(\U1761/U31/Z ), .e(
        \nchdr_ack[2] ), .f(\U1761/U31/Z ) );
    inv_1 \U1761/U31/U30/Uinv  ( .x(\U1761/U31/Z ), .a(\U1761/x[1] ) );
    aoi222_1 \U1632/U30/U1  ( .x(net178), .a(cack), .b(chdrctrlack), .c(cack), 
        .d(\U1632/Z ), .e(chdrctrlack), .f(\U1632/Z ) );
    inv_1 \U1632/U30/Uinv  ( .x(\U1632/Z ), .a(net178) );
    aoi222_1 \U1676/U30/U1  ( .x(hdrcd), .a(\chdrack[0] ), .b(\chdrack[1] ), 
        .c(\chdrack[0] ), .d(\U1676/Z ), .e(\chdrack[1] ), .f(\U1676/Z ) );
    inv_1 \U1676/U30/Uinv  ( .x(\U1676/Z ), .a(hdrcd) );
    nor3_1 \U1770/U21/Unr  ( .x(\U1770/U21/nr ), .a(\nchdr_ack[10] ), .b(
        \nchdr_ack[9] ), .c(\nchdr_ack[8] ) );
    nand3_1 \U1770/U21/Und  ( .x(\U1770/U21/nd ), .a(\nchdr_ack[10] ), .b(
        \nchdr_ack[9] ), .c(\nchdr_ack[8] ) );
    oa21_1 \U1770/U21/U1  ( .x(\U1770/U21/n2 ), .a(\U1770/U21/n2 ), .b(
        \U1770/U21/nr ), .c(\U1770/U21/nd ) );
    inv_1 \U1770/U21/U3  ( .x(\chdrack[1] ), .a(\U1770/U21/n2 ) );
    nor2_1 \U1652_0_/U2/U5  ( .x(\nchdr_ack[0] ), .a(\net242[10] ), .b(
        \net244[10] ) );
    ao222_2 \U1652_0_/U12/U19/U1/U1  ( .x(\net244[10] ), .a(\net243[10] ), .b(
        csize[0]), .c(\net243[10] ), .d(\net244[10] ), .e(csize[0]), .f(
        \net244[10] ) );
    ao222_2 \U1652_0_/U11/U19/U1/U1  ( .x(\net242[10] ), .a(csize[2]), .b(
        \net243[10] ), .c(csize[2]), .d(\net242[10] ), .e(\net243[10] ), .f(
        \net242[10] ) );
    nor2_1 \U1652_1_/U2/U5  ( .x(\nchdr_ack[1] ), .a(\net242[9] ), .b(
        \net244[9] ) );
    ao222_2 \U1652_1_/U12/U19/U1/U1  ( .x(\net244[9] ), .a(\net243[9] ), .b(
        csize[1]), .c(\net243[9] ), .d(\net244[9] ), .e(csize[1]), .f(
        \net244[9] ) );
    ao222_2 \U1652_1_/U11/U19/U1/U1  ( .x(\net242[9] ), .a(csize[3]), .b(
        \net243[9] ), .c(csize[3]), .d(\net242[9] ), .e(\net243[9] ), .f(
        \net242[9] ) );
    nor2_1 \U1652_2_/U2/U5  ( .x(\nchdr_ack[2] ), .a(\net242[8] ), .b(
        \net244[8] ) );
    ao222_2 \U1652_2_/U12/U19/U1/U1  ( .x(\net244[8] ), .a(\net243[8] ), .b(
        crnw[0]), .c(\net243[8] ), .d(\net244[8] ), .e(crnw[0]), .f(
        \net244[8] ) );
    ao222_2 \U1652_2_/U11/U19/U1/U1  ( .x(\net242[8] ), .a(crnw[1]), .b(
        \net243[8] ), .c(crnw[1]), .d(\net242[8] ), .e(\net243[8] ), .f(
        \net242[8] ) );
    nor2_1 \U1652_3_/U2/U5  ( .x(\nchdr_ack[3] ), .a(\net242[7] ), .b(
        \net244[7] ) );
    ao222_2 \U1652_3_/U12/U19/U1/U1  ( .x(\net244[7] ), .a(\net243[7] ), .b(
        ctag[0]), .c(\net243[7] ), .d(\net244[7] ), .e(ctag[0]), .f(
        \net244[7] ) );
    ao222_2 \U1652_3_/U11/U19/U1/U1  ( .x(\net242[7] ), .a(ctag[5]), .b(
        \net243[7] ), .c(ctag[5]), .d(\net242[7] ), .e(\net243[7] ), .f(
        \net242[7] ) );
    nor2_1 \U1652_4_/U2/U5  ( .x(\nchdr_ack[4] ), .a(\net242[6] ), .b(
        \net244[6] ) );
    ao222_2 \U1652_4_/U12/U19/U1/U1  ( .x(\net244[6] ), .a(\net243[6] ), .b(
        ctag[1]), .c(\net243[6] ), .d(\net244[6] ), .e(ctag[1]), .f(
        \net244[6] ) );
    ao222_2 \U1652_4_/U11/U19/U1/U1  ( .x(\net242[6] ), .a(ctag[6]), .b(
        \net243[6] ), .c(ctag[6]), .d(\net242[6] ), .e(\net243[6] ), .f(
        \net242[6] ) );
    nor2_1 \U1652_5_/U2/U5  ( .x(\nchdr_ack[5] ), .a(\net242[5] ), .b(
        \net244[5] ) );
    ao222_2 \U1652_5_/U12/U19/U1/U1  ( .x(\net244[5] ), .a(\net243[5] ), .b(
        ctag[2]), .c(\net243[5] ), .d(\net244[5] ), .e(ctag[2]), .f(
        \net244[5] ) );
    ao222_2 \U1652_5_/U11/U19/U1/U1  ( .x(\net242[5] ), .a(ctag[7]), .b(
        \net243[5] ), .c(ctag[7]), .d(\net242[5] ), .e(\net243[5] ), .f(
        \net242[5] ) );
    nor2_1 \U1652_6_/U2/U5  ( .x(\nchdr_ack[6] ), .a(\net242[4] ), .b(
        \net244[4] ) );
    ao222_2 \U1652_6_/U12/U19/U1/U1  ( .x(\net244[4] ), .a(\net243[4] ), .b(
        ctag[3]), .c(\net243[4] ), .d(\net244[4] ), .e(ctag[3]), .f(
        \net244[4] ) );
    ao222_2 \U1652_6_/U11/U19/U1/U1  ( .x(\net242[4] ), .a(ctag[8]), .b(
        \net243[4] ), .c(ctag[8]), .d(\net242[4] ), .e(\net243[4] ), .f(
        \net242[4] ) );
    nor2_1 \U1652_7_/U2/U5  ( .x(\nchdr_ack[7] ), .a(\net242[3] ), .b(
        \net244[3] ) );
    ao222_2 \U1652_7_/U12/U19/U1/U1  ( .x(\net244[3] ), .a(\net243[3] ), .b(
        ctag[4]), .c(\net243[3] ), .d(\net244[3] ), .e(ctag[4]), .f(
        \net244[3] ) );
    ao222_2 \U1652_7_/U11/U19/U1/U1  ( .x(\net242[3] ), .a(ctag[9]), .b(
        \net243[3] ), .c(ctag[9]), .d(\net242[3] ), .e(\net243[3] ), .f(
        \net242[3] ) );
    nor2_1 \U1652_8_/U2/U5  ( .x(\nchdr_ack[8] ), .a(\net242[2] ), .b(
        \net244[2] ) );
    ao222_2 \U1652_8_/U12/U19/U1/U1  ( .x(\net244[2] ), .a(\net243[2] ), .b(
        ccol[0]), .c(\net243[2] ), .d(\net244[2] ), .e(ccol[0]), .f(
        \net244[2] ) );
    ao222_2 \U1652_8_/U11/U19/U1/U1  ( .x(\net242[2] ), .a(ccol[3]), .b(
        \net243[2] ), .c(ccol[3]), .d(\net242[2] ), .e(\net243[2] ), .f(
        \net242[2] ) );
    nor2_1 \U1652_9_/U2/U5  ( .x(\nchdr_ack[9] ), .a(\net242[1] ), .b(
        \net244[1] ) );
    ao222_2 \U1652_9_/U12/U19/U1/U1  ( .x(\net244[1] ), .a(\net243[1] ), .b(
        ccol[1]), .c(\net243[1] ), .d(\net244[1] ), .e(ccol[1]), .f(
        \net244[1] ) );
    ao222_2 \U1652_9_/U11/U19/U1/U1  ( .x(\net242[1] ), .a(ccol[4]), .b(
        \net243[1] ), .c(ccol[4]), .d(\net242[1] ), .e(\net243[1] ), .f(
        \net242[1] ) );
    nor2_1 \U1652_10_/U2/U5  ( .x(\nchdr_ack[10] ), .a(\net242[0] ), .b(
        \net244[0] ) );
    ao222_2 \U1652_10_/U12/U19/U1/U1  ( .x(\net244[0] ), .a(\net243[0] ), .b(
        ccol[2]), .c(\net243[0] ), .d(\net244[0] ), .e(ccol[2]), .f(
        \net244[0] ) );
    ao222_2 \U1652_10_/U11/U19/U1/U1  ( .x(\net242[0] ), .a(ccol[5]), .b(
        \net243[0] ), .c(ccol[5]), .d(\net242[0] ), .e(\net243[0] ), .f(
        \net242[0] ) );
    nor2_1 \U1574_0_/U2/U5  ( .x(\U1574_0_/net231 ), .a(\rhdr_l[5] ), .b(
        \rhdr_h[5] ) );
    and2_1 \U1574_0_/U13/U8  ( .x(\net243[10] ), .a(\U1574_0_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_0_/U12/U19/U1/U1  ( .x(\rhdr_h[5] ), .a(n8), .b(
        \net242[10] ), .c(n8), .d(\rhdr_h[5] ), .e(\net242[10] ), .f(
        \rhdr_h[5] ) );
    ao222_2 \U1574_0_/U11/U19/U1/U1  ( .x(\rhdr_l[5] ), .a(\net244[10] ), .b(
        n7), .c(\net244[10] ), .d(\rhdr_l[5] ), .e(n8), .f(\rhdr_l[5] ) );
    nor2_1 \U1574_1_/U2/U5  ( .x(\U1574_1_/net231 ), .a(\rhdr_l[6] ), .b(
        \rhdr_h[6] ) );
    and2_1 \U1574_1_/U13/U8  ( .x(\net243[9] ), .a(\U1574_1_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_1_/U12/U19/U1/U1  ( .x(\rhdr_h[6] ), .a(n7), .b(\net242[9] 
        ), .c(n6), .d(\rhdr_h[6] ), .e(\net242[9] ), .f(\rhdr_h[6] ) );
    ao222_2 \U1574_1_/U11/U19/U1/U1  ( .x(\rhdr_l[6] ), .a(\net244[9] ), .b(n7
        ), .c(\net244[9] ), .d(\rhdr_l[6] ), .e(n8), .f(\rhdr_l[6] ) );
    nor2_1 \U1574_2_/U2/U5  ( .x(\U1574_2_/net231 ), .a(\rhdr_l[7] ), .b(
        \rhdr_h[7] ) );
    and2_1 \U1574_2_/U13/U8  ( .x(\net243[8] ), .a(\U1574_2_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_2_/U12/U19/U1/U1  ( .x(\rhdr_h[7] ), .a(n6), .b(\net242[8] 
        ), .c(n6), .d(\rhdr_h[7] ), .e(\net242[8] ), .f(\rhdr_h[7] ) );
    ao222_2 \U1574_2_/U11/U19/U1/U1  ( .x(\rhdr_l[7] ), .a(\net244[8] ), .b(n7
        ), .c(\net244[8] ), .d(\rhdr_l[7] ), .e(n8), .f(\rhdr_l[7] ) );
    nor2_1 \U1574_3_/U2/U5  ( .x(\U1574_3_/net231 ), .a(tag_l[0]), .b(tag_h[0]
        ) );
    and2_1 \U1574_3_/U13/U8  ( .x(\net243[7] ), .a(\U1574_3_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_3_/U12/U19/U1/U1  ( .x(tag_h[0]), .a(n8), .b(\net242[7] ), 
        .c(n6), .d(tag_h[0]), .e(\net242[7] ), .f(tag_h[0]) );
    ao222_2 \U1574_3_/U11/U19/U1/U1  ( .x(tag_l[0]), .a(\net244[7] ), .b(n7), 
        .c(\net244[7] ), .d(tag_l[0]), .e(n6), .f(tag_l[0]) );
    nor2_1 \U1574_4_/U2/U5  ( .x(\U1574_4_/net231 ), .a(tag_l[1]), .b(tag_h[1]
        ) );
    and2_1 \U1574_4_/U13/U8  ( .x(\net243[6] ), .a(\U1574_4_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_4_/U12/U19/U1/U1  ( .x(tag_h[1]), .a(n6), .b(\net242[6] ), 
        .c(n6), .d(tag_h[1]), .e(\net242[6] ), .f(tag_h[1]) );
    ao222_2 \U1574_4_/U11/U19/U1/U1  ( .x(tag_l[1]), .a(\net244[6] ), .b(n7), 
        .c(\net244[6] ), .d(tag_l[1]), .e(n6), .f(tag_l[1]) );
    nor2_1 \U1574_5_/U2/U5  ( .x(\U1574_5_/net231 ), .a(tag_l[2]), .b(tag_h[2]
        ) );
    and2_1 \U1574_5_/U13/U8  ( .x(\net243[5] ), .a(\U1574_5_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_5_/U12/U19/U1/U1  ( .x(tag_h[2]), .a(n7), .b(\net242[5] ), 
        .c(n6), .d(tag_h[2]), .e(\net242[5] ), .f(tag_h[2]) );
    ao222_2 \U1574_5_/U11/U19/U1/U1  ( .x(tag_l[2]), .a(\net244[5] ), .b(n7), 
        .c(\net244[5] ), .d(tag_l[2]), .e(n8), .f(tag_l[2]) );
    nor2_1 \U1574_6_/U2/U5  ( .x(\U1574_6_/net231 ), .a(tag_l[3]), .b(tag_h[3]
        ) );
    and2_1 \U1574_6_/U13/U8  ( .x(\net243[4] ), .a(\U1574_6_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_6_/U12/U19/U1/U1  ( .x(tag_h[3]), .a(n6), .b(\net242[4] ), 
        .c(n8), .d(tag_h[3]), .e(\net242[4] ), .f(tag_h[3]) );
    ao222_2 \U1574_6_/U11/U19/U1/U1  ( .x(tag_l[3]), .a(\net244[4] ), .b(n7), 
        .c(\net244[4] ), .d(tag_l[3]), .e(n6), .f(tag_l[3]) );
    nor2_1 \U1574_7_/U2/U5  ( .x(\U1574_7_/net231 ), .a(tag_l[4]), .b(tag_h[4]
        ) );
    and2_1 \U1574_7_/U13/U8  ( .x(\net243[3] ), .a(\U1574_7_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_7_/U12/U19/U1/U1  ( .x(tag_h[4]), .a(n6), .b(\net242[3] ), 
        .c(n8), .d(tag_h[4]), .e(\net242[3] ), .f(tag_h[4]) );
    ao222_2 \U1574_7_/U11/U19/U1/U1  ( .x(tag_l[4]), .a(\net244[3] ), .b(n7), 
        .c(\net244[3] ), .d(tag_l[4]), .e(n6), .f(tag_l[4]) );
    nor2_1 \U1574_8_/U2/U5  ( .x(\U1574_8_/net231 ), .a(\rhdr_l[13] ), .b(
        \rhdr_h[13] ) );
    and2_1 \U1574_8_/U13/U8  ( .x(\net243[2] ), .a(\U1574_8_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_8_/U12/U19/U1/U1  ( .x(\rhdr_h[13] ), .a(n7), .b(
        \net242[2] ), .c(n8), .d(\rhdr_h[13] ), .e(\net242[2] ), .f(
        \rhdr_h[13] ) );
    ao222_2 \U1574_8_/U11/U19/U1/U1  ( .x(\rhdr_l[13] ), .a(\net244[2] ), .b(
        n7), .c(\net244[2] ), .d(\rhdr_l[13] ), .e(n6), .f(\rhdr_l[13] ) );
    nor2_1 \U1574_9_/U2/U5  ( .x(\U1574_9_/net231 ), .a(\rhdr_l[14] ), .b(
        \rhdr_h[14] ) );
    and2_1 \U1574_9_/U13/U8  ( .x(\net243[1] ), .a(\U1574_9_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_9_/U12/U19/U1/U1  ( .x(\rhdr_h[14] ), .a(n8), .b(
        \net242[1] ), .c(n6), .d(\rhdr_h[14] ), .e(\net242[1] ), .f(
        \rhdr_h[14] ) );
    ao222_2 \U1574_9_/U11/U19/U1/U1  ( .x(\rhdr_l[14] ), .a(\net244[1] ), .b(
        n7), .c(\net244[1] ), .d(\rhdr_l[14] ), .e(n8), .f(\rhdr_l[14] ) );
    nor2_1 \U1574_10_/U2/U5  ( .x(\U1574_10_/net231 ), .a(\rhdr_l[15] ), .b(
        \rhdr_h[15] ) );
    and2_1 \U1574_10_/U13/U8  ( .x(\net243[0] ), .a(\U1574_10_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_10_/U12/U19/U1/U1  ( .x(\rhdr_h[15] ), .a(n8), .b(
        \net242[0] ), .c(n8), .d(\rhdr_h[15] ), .e(\net242[0] ), .f(
        \rhdr_h[15] ) );
    ao222_2 \U1574_10_/U11/U19/U1/U1  ( .x(\rhdr_l[15] ), .a(\net244[0] ), .b(
        n7), .c(\net244[0] ), .d(\rhdr_l[15] ), .e(n8), .f(\rhdr_l[15] ) );
    buf_1 U1 ( .x(csize[0]), .a(n12) );
    buf_1 U2 ( .x(csize[1]), .a(n11) );
    buf_1 U3 ( .x(crnw[0]), .a(n10) );
    buf_1 U4 ( .x(crnw[1]), .a(n9) );
    inv_5 U5 ( .x(n5), .a(net265) );
    buf_3 U6 ( .x(nbreset), .a(nReset) );
    buf_3 U7 ( .x(n6), .a(net248) );
    buf_3 U8 ( .x(n8), .a(net248) );
    buf_3 U9 ( .x(n7), .a(net248) );
    nor2_1 U10 ( .x(net248), .a(net265), .b(rhdrack) );
endmodule


module chain_selement_ga_16 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_15 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[1] , \c[0] ;
    chain_selement_ga_16 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_17 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_16 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[1] , \c[0] ;
    chain_selement_ga_17 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_18 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_17 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[1] , \c[0] , n1, n2;
    chain_selement_ga_18 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        n2), .e(n2) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(n2), .b(r[0]), .c(n2), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(n2), .b(r[1]), .c(n2), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
    inv_0 U1 ( .x(n1), .a(e[0]) );
    inv_2 U2 ( .x(n2), .a(n1) );
endmodule


module chain_selement_ga_75 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module resp_route_tx_imem ( o, rtxack, e_h, e_l, noa, r_h, r_l, rtxreq );
output [4:0] o;
input  [2:0] e_h;
input  [2:0] e_l;
input  [2:0] r_h;
input  [2:0] r_l;
input  noa, rtxreq;
output rtxack;
    wire \r2[2] , \r2[1] , \r2[0] , \r1[2] , \r1[1] , \r1[0] , \r0[2] , 
        \r0[1] , \r0[0] , \last[0] , \last[1] , \last[2] , \last[3] , 
        \net72[0] , \net72[1] , net56, net106, net103, eopsym, net87, net66, 
        net84, net77, \I8/nb , \I8/na , \I11/n5 , \I11/n1 , \I11/n2 , \I11/n3 , 
        \I11/n4 , \I7_0_/U25/U1/clr , \I7_0_/U25/U1/ob , \I7_1_/U25/U1/clr , 
        \I7_1_/U25/U1/ob ;
    assign o[3] = 1'b0;
    assign o[2] = 1'b0;
    chain_selement_ga_75 I9 ( .Aa(\last[0] ), .Br(eopsym), .Ar(net87), .Ba(
        net66) );
    route_symbol_16 I2 ( .o({\r1[2] , \r1[1] , \r1[0] }), .txack(net84), 
        .txack_last(\last[2] ), .e({e_h[1], e_l[1]}), .oa(net66), .r({r_h[1], 
        r_l[1]}), .txreq(net77) );
    route_symbol_17 I3 ( .o({\r0[2] , \r0[1] , \r0[0] }), .txack(net87), 
        .txack_last(\last[1] ), .e({e_h[0], e_l[0]}), .oa(net66), .r({r_h[0], 
        r_l[0]}), .txreq(net84) );
    route_symbol_15 I1 ( .o({\r2[2] , \r2[1] , \r2[0] }), .txack(net77), 
        .txack_last(\last[3] ), .e({e_h[2], e_l[2]}), .oa(net66), .r({r_h[2], 
        r_l[2]}), .txreq(rtxreq) );
    nor2_1 \I5/U5  ( .x(net106), .a(eopsym), .b(\r2[2] ) );
    nor2_1 \I16/U5  ( .x(net103), .a(\r1[2] ), .b(\r0[2] ) );
    or2_1 \I14_0_/U12  ( .x(\net72[1] ), .a(\r2[0] ), .b(\r1[0] ) );
    or2_1 \I14_1_/U12  ( .x(\net72[0] ), .a(\r2[1] ), .b(\r1[1] ) );
    nor3_1 \I8/U27  ( .x(\I8/nb ), .a(o[4]), .b(o[3]), .c(o[2]) );
    nor2_1 \I8/U26  ( .x(\I8/na ), .a(o[1]), .b(o[0]) );
    nand2_2 \I8/U29  ( .x(net66), .a(\I8/nb ), .b(\I8/na ) );
    and4_1 \I11/U16  ( .x(\I11/n5 ), .a(\I11/n1 ), .b(\I11/n2 ), .c(\I11/n3 ), 
        .d(\I11/n4 ) );
    inv_1 \I11/U1  ( .x(\I11/n1 ), .a(\last[3] ) );
    inv_1 \I11/U2  ( .x(\I11/n2 ), .a(\last[2] ) );
    inv_1 \I11/U3  ( .x(\I11/n3 ), .a(\last[1] ) );
    inv_1 \I11/U4  ( .x(\I11/n4 ), .a(\last[0] ) );
    inv_1 \I11/U5  ( .x(rtxack), .a(\I11/n5 ) );
    nand2_1 \I17/U5  ( .x(net56), .a(net106), .b(net103) );
    ao222_1 \I15/U18/U1/U1  ( .x(o[4]), .a(noa), .b(net56), .c(noa), .d(o[4]), 
        .e(net56), .f(o[4]) );
    oa31_1 \I7_0_/U25/U1/Uclr  ( .x(\I7_0_/U25/U1/clr ), .a(noa), .b(\r0[0] ), 
        .c(\net72[1] ), .d(o[0]) );
    oaoi211_1 \I7_0_/U25/U1/Uaoi  ( .x(\I7_0_/U25/U1/ob ), .a(\r0[0] ), .b(
        \net72[1] ), .c(noa), .d(\I7_0_/U25/U1/clr ) );
    inv_2 \I7_0_/U25/U1/Ui  ( .x(o[0]), .a(\I7_0_/U25/U1/ob ) );
    oa31_1 \I7_1_/U25/U1/Uclr  ( .x(\I7_1_/U25/U1/clr ), .a(noa), .b(\r0[1] ), 
        .c(\net72[0] ), .d(o[1]) );
    oaoi211_1 \I7_1_/U25/U1/Uaoi  ( .x(\I7_1_/U25/U1/ob ), .a(\r0[1] ), .b(
        \net72[0] ), .c(noa), .d(\I7_1_/U25/U1/clr ) );
    inv_2 \I7_1_/U25/U1/Ui  ( .x(o[1]), .a(\I7_1_/U25/U1/ob ) );
endmodule


module matched_delay_cp2slave_resp_imem ( x, a );
input  a;
output x;
    buf_1 I1 ( .x(x), .a(a) );
endmodule


module matched_delay_cp2slave_comimem ( x, a );
input  a;
output x;
    buf_1 I1 ( .x(x), .a(a) );
endmodule


module sr2dr_word_7 ( i, req, h, l );
input  [31:0] i;
output [31:0] h;
output [31:0] l;
input  req;
    wire \U31/nl , \U31/ni , \U31/nh , \U30/nl , \U30/ni , \U30/nh , \U29/nl , 
        \U29/ni , \U29/nh , \U28/nl , \U28/ni , \U28/nh , \U27/nl , \U27/ni , 
        \U27/nh , \U26/nl , \U26/ni , \U26/nh , \U25/nl , \U25/ni , \U25/nh , 
        \U24/nl , \U24/ni , \U24/nh , \U23/nl , \U23/ni , \U23/nh , \U22/nl , 
        \U22/ni , \U22/nh , \U21/nl , \U21/ni , \U21/nh , \U20/nl , \U20/ni , 
        \U20/nh , \U19/nl , \U19/ni , \U19/nh , \U18/nl , \U18/ni , \U18/nh , 
        \U17/nl , \U17/ni , \U17/nh , \U16/nl , \U16/ni , \U16/nh , \U15/nl , 
        \U15/ni , \U15/nh , \U14/nl , \U14/ni , \U14/nh , \U13/nl , \U13/ni , 
        \U13/nh , \U12/nl , \U12/ni , \U12/nh , \U11/nl , \U11/ni , \U11/nh , 
        \U10/nl , \U10/ni , \U10/nh , \U9/nl , \U9/ni , \U9/nh , \U8/nl , 
        \U8/ni , \U8/nh , \U7/nl , \U7/ni , \U7/nh , \U6/nl , \U6/ni , \U6/nh , 
        \U5/nl , \U5/ni , \U5/nh , \U4/nl , \U4/ni , \U4/nh , \U3/nl , \U3/ni , 
        \U3/nh , \U2/nl , \U2/ni , \U2/nh , \U1/nl , \U1/ni , \U1/nh , \U0/nl , 
        \U0/ni , \U0/nh , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
    inv_1 \U31/Uii  ( .x(\U31/ni ), .a(i[31]) );
    inv_1 \U31/Uih  ( .x(\U31/nh ), .a(h[31]) );
    inv_1 \U31/Uil  ( .x(\U31/nl ), .a(l[31]) );
    ao23_1 \U31/Ucl/U1/U1  ( .x(l[31]), .a(n9), .b(l[31]), .c(n1), .d(\U31/ni 
        ), .e(\U31/nh ) );
    ao23_1 \U31/Uch/U1/U1  ( .x(h[31]), .a(n9), .b(h[31]), .c(n2), .d(i[31]), 
        .e(\U31/nl ) );
    inv_1 \U30/Uii  ( .x(\U30/ni ), .a(i[30]) );
    inv_1 \U30/Uih  ( .x(\U30/nh ), .a(h[30]) );
    inv_1 \U30/Uil  ( .x(\U30/nl ), .a(l[30]) );
    ao23_1 \U30/Ucl/U1/U1  ( .x(l[30]), .a(n8), .b(l[30]), .c(n1), .d(\U30/ni 
        ), .e(\U30/nh ) );
    ao23_1 \U30/Uch/U1/U1  ( .x(h[30]), .a(n8), .b(h[30]), .c(n1), .d(i[30]), 
        .e(\U30/nl ) );
    inv_1 \U29/Uii  ( .x(\U29/ni ), .a(i[29]) );
    inv_1 \U29/Uih  ( .x(\U29/nh ), .a(h[29]) );
    inv_1 \U29/Uil  ( .x(\U29/nl ), .a(l[29]) );
    ao23_1 \U29/Ucl/U1/U1  ( .x(l[29]), .a(n8), .b(l[29]), .c(n1), .d(\U29/ni 
        ), .e(\U29/nh ) );
    ao23_1 \U29/Uch/U1/U1  ( .x(h[29]), .a(n8), .b(h[29]), .c(n2), .d(i[29]), 
        .e(\U29/nl ) );
    inv_1 \U28/Uii  ( .x(\U28/ni ), .a(i[28]) );
    inv_1 \U28/Uih  ( .x(\U28/nh ), .a(h[28]) );
    inv_1 \U28/Uil  ( .x(\U28/nl ), .a(l[28]) );
    ao23_1 \U28/Ucl/U1/U1  ( .x(l[28]), .a(n8), .b(l[28]), .c(n2), .d(\U28/ni 
        ), .e(\U28/nh ) );
    ao23_1 \U28/Uch/U1/U1  ( .x(h[28]), .a(n8), .b(h[28]), .c(n2), .d(i[28]), 
        .e(\U28/nl ) );
    inv_1 \U27/Uii  ( .x(\U27/ni ), .a(i[27]) );
    inv_1 \U27/Uih  ( .x(\U27/nh ), .a(h[27]) );
    inv_1 \U27/Uil  ( .x(\U27/nl ), .a(l[27]) );
    ao23_1 \U27/Ucl/U1/U1  ( .x(l[27]), .a(n8), .b(l[27]), .c(n2), .d(\U27/ni 
        ), .e(\U27/nh ) );
    ao23_1 \U27/Uch/U1/U1  ( .x(h[27]), .a(n8), .b(h[27]), .c(n2), .d(i[27]), 
        .e(\U27/nl ) );
    inv_1 \U26/Uii  ( .x(\U26/ni ), .a(i[26]) );
    inv_1 \U26/Uih  ( .x(\U26/nh ), .a(h[26]) );
    inv_1 \U26/Uil  ( .x(\U26/nl ), .a(l[26]) );
    ao23_1 \U26/Ucl/U1/U1  ( .x(l[26]), .a(n7), .b(l[26]), .c(n2), .d(\U26/ni 
        ), .e(\U26/nh ) );
    ao23_1 \U26/Uch/U1/U1  ( .x(h[26]), .a(n7), .b(h[26]), .c(n4), .d(i[26]), 
        .e(\U26/nl ) );
    inv_1 \U25/Uii  ( .x(\U25/ni ), .a(i[25]) );
    inv_1 \U25/Uih  ( .x(\U25/nh ), .a(h[25]) );
    inv_1 \U25/Uil  ( .x(\U25/nl ), .a(l[25]) );
    ao23_1 \U25/Ucl/U1/U1  ( .x(l[25]), .a(n7), .b(l[25]), .c(n4), .d(\U25/ni 
        ), .e(\U25/nh ) );
    ao23_1 \U25/Uch/U1/U1  ( .x(h[25]), .a(n7), .b(h[25]), .c(n4), .d(i[25]), 
        .e(\U25/nl ) );
    inv_1 \U24/Uii  ( .x(\U24/ni ), .a(i[24]) );
    inv_1 \U24/Uih  ( .x(\U24/nh ), .a(h[24]) );
    inv_1 \U24/Uil  ( .x(\U24/nl ), .a(l[24]) );
    ao23_1 \U24/Ucl/U1/U1  ( .x(l[24]), .a(n7), .b(l[24]), .c(n4), .d(\U24/ni 
        ), .e(\U24/nh ) );
    ao23_1 \U24/Uch/U1/U1  ( .x(h[24]), .a(n7), .b(h[24]), .c(n4), .d(i[24]), 
        .e(\U24/nl ) );
    inv_1 \U23/Uii  ( .x(\U23/ni ), .a(i[23]) );
    inv_1 \U23/Uih  ( .x(\U23/nh ), .a(h[23]) );
    inv_1 \U23/Uil  ( .x(\U23/nl ), .a(l[23]) );
    ao23_1 \U23/Ucl/U1/U1  ( .x(l[23]), .a(n7), .b(l[23]), .c(n3), .d(\U23/ni 
        ), .e(\U23/nh ) );
    ao23_1 \U23/Uch/U1/U1  ( .x(h[23]), .a(n7), .b(h[23]), .c(n3), .d(i[23]), 
        .e(\U23/nl ) );
    inv_1 \U22/Uii  ( .x(\U22/ni ), .a(i[22]) );
    inv_1 \U22/Uih  ( .x(\U22/nh ), .a(h[22]) );
    inv_1 \U22/Uil  ( .x(\U22/nl ), .a(l[22]) );
    ao23_1 \U22/Ucl/U1/U1  ( .x(l[22]), .a(n6), .b(l[22]), .c(n3), .d(\U22/ni 
        ), .e(\U22/nh ) );
    ao23_1 \U22/Uch/U1/U1  ( .x(h[22]), .a(n6), .b(h[22]), .c(n3), .d(i[22]), 
        .e(\U22/nl ) );
    inv_1 \U21/Uii  ( .x(\U21/ni ), .a(i[21]) );
    inv_1 \U21/Uih  ( .x(\U21/nh ), .a(h[21]) );
    inv_1 \U21/Uil  ( .x(\U21/nl ), .a(l[21]) );
    ao23_1 \U21/Ucl/U1/U1  ( .x(l[21]), .a(n6), .b(l[21]), .c(n3), .d(\U21/ni 
        ), .e(\U21/nh ) );
    ao23_1 \U21/Uch/U1/U1  ( .x(h[21]), .a(n6), .b(h[21]), .c(n3), .d(i[21]), 
        .e(\U21/nl ) );
    inv_1 \U20/Uii  ( .x(\U20/ni ), .a(i[20]) );
    inv_1 \U20/Uih  ( .x(\U20/nh ), .a(h[20]) );
    inv_1 \U20/Uil  ( .x(\U20/nl ), .a(l[20]) );
    ao23_1 \U20/Ucl/U1/U1  ( .x(l[20]), .a(n6), .b(l[20]), .c(n5), .d(\U20/ni 
        ), .e(\U20/nh ) );
    ao23_1 \U20/Uch/U1/U1  ( .x(h[20]), .a(n6), .b(h[20]), .c(n4), .d(i[20]), 
        .e(\U20/nl ) );
    inv_1 \U19/Uii  ( .x(\U19/ni ), .a(i[19]) );
    inv_1 \U19/Uih  ( .x(\U19/nh ), .a(h[19]) );
    inv_1 \U19/Uil  ( .x(\U19/nl ), .a(l[19]) );
    ao23_1 \U19/Ucl/U1/U1  ( .x(l[19]), .a(n6), .b(l[19]), .c(n4), .d(\U19/ni 
        ), .e(\U19/nh ) );
    ao23_1 \U19/Uch/U1/U1  ( .x(h[19]), .a(n6), .b(h[19]), .c(n4), .d(i[19]), 
        .e(\U19/nl ) );
    inv_1 \U18/Uii  ( .x(\U18/ni ), .a(i[18]) );
    inv_1 \U18/Uih  ( .x(\U18/nh ), .a(h[18]) );
    inv_1 \U18/Uil  ( .x(\U18/nl ), .a(l[18]) );
    ao23_1 \U18/Ucl/U1/U1  ( .x(l[18]), .a(n5), .b(l[18]), .c(n5), .d(\U18/ni 
        ), .e(\U18/nh ) );
    ao23_1 \U18/Uch/U1/U1  ( .x(h[18]), .a(n5), .b(h[18]), .c(n5), .d(i[18]), 
        .e(\U18/nl ) );
    inv_1 \U17/Uii  ( .x(\U17/ni ), .a(i[17]) );
    inv_1 \U17/Uih  ( .x(\U17/nh ), .a(h[17]) );
    inv_1 \U17/Uil  ( .x(\U17/nl ), .a(l[17]) );
    ao23_1 \U17/Ucl/U1/U1  ( .x(l[17]), .a(n6), .b(l[17]), .c(n5), .d(\U17/ni 
        ), .e(\U17/nh ) );
    ao23_1 \U17/Uch/U1/U1  ( .x(h[17]), .a(n7), .b(h[17]), .c(n4), .d(i[17]), 
        .e(\U17/nl ) );
    inv_1 \U16/Uii  ( .x(\U16/ni ), .a(i[16]) );
    inv_1 \U16/Uih  ( .x(\U16/nh ), .a(h[16]) );
    inv_1 \U16/Uil  ( .x(\U16/nl ), .a(l[16]) );
    ao23_1 \U16/Ucl/U1/U1  ( .x(l[16]), .a(n9), .b(l[16]), .c(n3), .d(\U16/ni 
        ), .e(\U16/nh ) );
    ao23_1 \U16/Uch/U1/U1  ( .x(h[16]), .a(n9), .b(h[16]), .c(n1), .d(i[16]), 
        .e(\U16/nl ) );
    inv_1 \U15/Uii  ( .x(\U15/ni ), .a(i[15]) );
    inv_1 \U15/Uih  ( .x(\U15/nh ), .a(h[15]) );
    inv_1 \U15/Uil  ( .x(\U15/nl ), .a(l[15]) );
    ao23_1 \U15/Ucl/U1/U1  ( .x(l[15]), .a(n8), .b(l[15]), .c(n1), .d(\U15/ni 
        ), .e(\U15/nh ) );
    ao23_1 \U15/Uch/U1/U1  ( .x(h[15]), .a(n7), .b(h[15]), .c(n1), .d(i[15]), 
        .e(\U15/nl ) );
    inv_1 \U14/Uii  ( .x(\U14/ni ), .a(i[14]) );
    inv_1 \U14/Uih  ( .x(\U14/nh ), .a(h[14]) );
    inv_1 \U14/Uil  ( .x(\U14/nl ), .a(l[14]) );
    ao23_1 \U14/Ucl/U1/U1  ( .x(l[14]), .a(n6), .b(l[14]), .c(n1), .d(\U14/ni 
        ), .e(\U14/nh ) );
    ao23_1 \U14/Uch/U1/U1  ( .x(h[14]), .a(n6), .b(h[14]), .c(n3), .d(i[14]), 
        .e(\U14/nl ) );
    inv_1 \U13/Uii  ( .x(\U13/ni ), .a(i[13]) );
    inv_1 \U13/Uih  ( .x(\U13/nh ), .a(h[13]) );
    inv_1 \U13/Uil  ( .x(\U13/nl ), .a(l[13]) );
    ao23_1 \U13/Ucl/U1/U1  ( .x(l[13]), .a(n6), .b(l[13]), .c(n4), .d(\U13/ni 
        ), .e(\U13/nh ) );
    ao23_1 \U13/Uch/U1/U1  ( .x(h[13]), .a(n6), .b(h[13]), .c(n4), .d(i[13]), 
        .e(\U13/nl ) );
    inv_1 \U12/Uii  ( .x(\U12/ni ), .a(i[12]) );
    inv_1 \U12/Uih  ( .x(\U12/nh ), .a(h[12]) );
    inv_1 \U12/Uil  ( .x(\U12/nl ), .a(l[12]) );
    ao23_1 \U12/Ucl/U1/U1  ( .x(l[12]), .a(n5), .b(l[12]), .c(n4), .d(\U12/ni 
        ), .e(\U12/nh ) );
    ao23_1 \U12/Uch/U1/U1  ( .x(h[12]), .a(n5), .b(h[12]), .c(n4), .d(i[12]), 
        .e(\U12/nl ) );
    inv_1 \U11/Uii  ( .x(\U11/ni ), .a(i[11]) );
    inv_1 \U11/Uih  ( .x(\U11/nh ), .a(h[11]) );
    inv_1 \U11/Uil  ( .x(\U11/nl ), .a(l[11]) );
    ao23_1 \U11/Ucl/U1/U1  ( .x(l[11]), .a(n5), .b(l[11]), .c(n4), .d(\U11/ni 
        ), .e(\U11/nh ) );
    ao23_1 \U11/Uch/U1/U1  ( .x(h[11]), .a(n5), .b(h[11]), .c(n4), .d(i[11]), 
        .e(\U11/nl ) );
    inv_1 \U10/Uii  ( .x(\U10/ni ), .a(i[10]) );
    inv_1 \U10/Uih  ( .x(\U10/nh ), .a(h[10]) );
    inv_1 \U10/Uil  ( .x(\U10/nl ), .a(l[10]) );
    ao23_1 \U10/Ucl/U1/U1  ( .x(l[10]), .a(n5), .b(l[10]), .c(n3), .d(\U10/ni 
        ), .e(\U10/nh ) );
    ao23_1 \U10/Uch/U1/U1  ( .x(h[10]), .a(n5), .b(h[10]), .c(n3), .d(i[10]), 
        .e(\U10/nl ) );
    inv_1 \U9/Uii  ( .x(\U9/ni ), .a(i[9]) );
    inv_1 \U9/Uih  ( .x(\U9/nh ), .a(h[9]) );
    inv_1 \U9/Uil  ( .x(\U9/nl ), .a(l[9]) );
    ao23_1 \U9/Ucl/U1/U1  ( .x(l[9]), .a(n5), .b(l[9]), .c(n3), .d(\U9/ni ), 
        .e(\U9/nh ) );
    ao23_1 \U9/Uch/U1/U1  ( .x(h[9]), .a(n5), .b(h[9]), .c(n3), .d(i[9]), .e(
        \U9/nl ) );
    inv_1 \U8/Uii  ( .x(\U8/ni ), .a(i[8]) );
    inv_1 \U8/Uih  ( .x(\U8/nh ), .a(h[8]) );
    inv_1 \U8/Uil  ( .x(\U8/nl ), .a(l[8]) );
    ao23_1 \U8/Ucl/U1/U1  ( .x(l[8]), .a(n5), .b(l[8]), .c(n3), .d(\U8/ni ), 
        .e(\U8/nh ) );
    ao23_1 \U8/Uch/U1/U1  ( .x(h[8]), .a(n5), .b(h[8]), .c(n3), .d(i[8]), .e(
        \U8/nl ) );
    inv_1 \U7/Uii  ( .x(\U7/ni ), .a(i[7]) );
    inv_1 \U7/Uih  ( .x(\U7/nh ), .a(h[7]) );
    inv_1 \U7/Uil  ( .x(\U7/nl ), .a(l[7]) );
    ao23_1 \U7/Ucl/U1/U1  ( .x(l[7]), .a(n7), .b(l[7]), .c(n3), .d(\U7/ni ), 
        .e(\U7/nh ) );
    ao23_1 \U7/Uch/U1/U1  ( .x(h[7]), .a(n7), .b(h[7]), .c(n2), .d(i[7]), .e(
        \U7/nl ) );
    inv_1 \U6/Uii  ( .x(\U6/ni ), .a(i[6]) );
    inv_1 \U6/Uih  ( .x(\U6/nh ), .a(h[6]) );
    inv_1 \U6/Uil  ( .x(\U6/nl ), .a(l[6]) );
    ao23_1 \U6/Ucl/U1/U1  ( .x(l[6]), .a(n7), .b(l[6]), .c(n2), .d(\U6/ni ), 
        .e(\U6/nh ) );
    ao23_1 \U6/Uch/U1/U1  ( .x(h[6]), .a(n7), .b(h[6]), .c(n2), .d(i[6]), .e(
        \U6/nl ) );
    inv_1 \U5/Uii  ( .x(\U5/ni ), .a(i[5]) );
    inv_1 \U5/Uih  ( .x(\U5/nh ), .a(h[5]) );
    inv_1 \U5/Uil  ( .x(\U5/nl ), .a(l[5]) );
    ao23_1 \U5/Ucl/U1/U1  ( .x(l[5]), .a(n7), .b(l[5]), .c(n2), .d(\U5/ni ), 
        .e(\U5/nh ) );
    ao23_1 \U5/Uch/U1/U1  ( .x(h[5]), .a(n7), .b(h[5]), .c(n2), .d(i[5]), .e(
        \U5/nl ) );
    inv_1 \U4/Uii  ( .x(\U4/ni ), .a(i[4]) );
    inv_1 \U4/Uih  ( .x(\U4/nh ), .a(h[4]) );
    inv_1 \U4/Uil  ( .x(\U4/nl ), .a(l[4]) );
    ao23_1 \U4/Ucl/U1/U1  ( .x(l[4]), .a(n6), .b(l[4]), .c(n2), .d(\U4/ni ), 
        .e(\U4/nh ) );
    ao23_1 \U4/Uch/U1/U1  ( .x(h[4]), .a(n6), .b(h[4]), .c(n2), .d(i[4]), .e(
        \U4/nl ) );
    inv_1 \U3/Uii  ( .x(\U3/ni ), .a(i[3]) );
    inv_1 \U3/Uih  ( .x(\U3/nh ), .a(h[3]) );
    inv_1 \U3/Uil  ( .x(\U3/nl ), .a(l[3]) );
    ao23_1 \U3/Ucl/U1/U1  ( .x(l[3]), .a(n6), .b(l[3]), .c(n2), .d(\U3/ni ), 
        .e(\U3/nh ) );
    ao23_1 \U3/Uch/U1/U1  ( .x(h[3]), .a(n8), .b(h[3]), .c(n1), .d(i[3]), .e(
        \U3/nl ) );
    inv_1 \U2/Uii  ( .x(\U2/ni ), .a(i[2]) );
    inv_1 \U2/Uih  ( .x(\U2/nh ), .a(h[2]) );
    inv_1 \U2/Uil  ( .x(\U2/nl ), .a(l[2]) );
    ao23_1 \U2/Ucl/U1/U1  ( .x(l[2]), .a(n8), .b(l[2]), .c(n1), .d(\U2/ni ), 
        .e(\U2/nh ) );
    ao23_1 \U2/Uch/U1/U1  ( .x(h[2]), .a(n8), .b(h[2]), .c(n1), .d(i[2]), .e(
        \U2/nl ) );
    inv_1 \U1/Uii  ( .x(\U1/ni ), .a(i[1]) );
    inv_1 \U1/Uih  ( .x(\U1/nh ), .a(h[1]) );
    inv_1 \U1/Uil  ( .x(\U1/nl ), .a(l[1]) );
    ao23_1 \U1/Ucl/U1/U1  ( .x(l[1]), .a(n8), .b(l[1]), .c(n1), .d(\U1/ni ), 
        .e(\U1/nh ) );
    ao23_1 \U1/Uch/U1/U1  ( .x(h[1]), .a(n8), .b(h[1]), .c(n1), .d(i[1]), .e(
        \U1/nl ) );
    inv_1 \U0/Uii  ( .x(\U0/ni ), .a(i[0]) );
    inv_1 \U0/Uih  ( .x(\U0/nh ), .a(h[0]) );
    inv_1 \U0/Uil  ( .x(\U0/nl ), .a(l[0]) );
    ao23_1 \U0/Ucl/U1/U1  ( .x(l[0]), .a(n8), .b(l[0]), .c(n1), .d(\U0/ni ), 
        .e(\U0/nh ) );
    ao23_1 \U0/Uch/U1/U1  ( .x(h[0]), .a(n8), .b(h[0]), .c(n1), .d(i[0]), .e(
        \U0/nl ) );
    buf_16 U1 ( .x(n1), .a(n12) );
    buf_16 U2 ( .x(n2), .a(n12) );
    buf_16 U3 ( .x(n3), .a(n12) );
    buf_16 U4 ( .x(n4), .a(n11) );
    buf_16 U5 ( .x(n5), .a(n11) );
    buf_16 U6 ( .x(n6), .a(n11) );
    buf_16 U7 ( .x(n7), .a(n10) );
    buf_16 U8 ( .x(n8), .a(n10) );
    buf_16 U9 ( .x(n9), .a(n10) );
    buf_16 U10 ( .x(n10), .a(req) );
    buf_16 U11 ( .x(n11), .a(req) );
    buf_16 U12 ( .x(n12), .a(req) );
endmodule


module cp2slave_imem ( tc_seq, tc_size, tc_itag, tc_wd, tc_lock, tc_a, tc_rnw, 
    tc_ok, tc_defer, tc_slow, tc_ack, req_in, ts_i, st_i, we_i, mult_i, adr_i, 
    dat_i, seq_i, prd_i, sel_i, ack_in, tr_rd, tr_err, tr_size, tr_ack, tr_rnw, 
    req_out, dat_o, err_o, rty_o, acc_o, sel_o, mult_o, rt_o, ack_out, reset
     );
input  [1:0] tc_seq;
input  [3:0] tc_size;
input  [9:0] tc_itag;
input  [63:0] tc_wd;
input  [1:0] tc_lock;
input  [63:0] tc_a;
input  [1:0] tc_rnw;
output [2:0] ts_i;
output [4:0] st_i;
output [31:0] adr_i;
output [31:0] dat_i;
output [3:0] sel_i;
output [63:0] tr_rd;
output [1:0] tr_err;
output [3:0] tr_size;
output [1:0] tr_rnw;
input  [31:0] dat_o;
input  [3:0] sel_o;
input  [4:0] rt_o;
input  ack_in, tr_ack, req_out, err_o, rty_o, acc_o, mult_o, reset;
output tc_ok, tc_defer, tc_slow, tc_ack, req_in, we_i, mult_i, seq_i, prd_i, 
    ack_out;
    wire \tc_a[60] , \tc_a[58] , \tc_wd[63] , \tc_wd[62] , \tc_wd[61] , 
        \tc_wd[60] , \tc_wd[59] , \tc_wd[58] , \tc_wd[56] , \tc_wd[55] , 
        \tc_wd[54] , \tc_wd[53] , \tc_wd[52] , \tc_wd[51] , \tc_wd[50] , 
        \tc_wd[49] , \tc_wd[48] , \tc_wd[47] , \tc_wd[46] , \tc_wd[45] , 
        \tc_wd[44] , \tc_wd[43] , \tc_wd[40] , \tc_wd[39] , \tc_wd[38] , 
        \tc_wd[36] , \tc_wd[32] , \sel_i[2] , n121, n122, n123, n124, n125, 
        n126, n127, n128, n129, n130, n135, n136, n137, n141, n142, n180, n181, 
        n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, 
        n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, 
        n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, 
        n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
        n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, 
        n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, 
        n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, 
        n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, 
        n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, 
        n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, 
        n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, 
        n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, 
        n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, 
        n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, 
        n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, 
        n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, 
        n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, 
        n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, 
        n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
        n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
        n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
        n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
        n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
        n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
        n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
        n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
        n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
        n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
        n518, n519, n520, n521, n522, n523, n524, n525, n529, n530, n531, n532, 
        n3, n4, n5, complb1, complb0, comp_basic, complw1, complw0, comp_wd, 
        all_w, all_r, respond, _24_net_, _25_net_, _26_net_, req_out_delayed, 
        req_in_i, \cg_all_w/__tmp99/loop , \Usze1/nl , \Usze1/ni , \Usze1/nh , 
        \Usze0/nl , \Usze0/ni , \Usze0/nh , \Urnw/nl , \Urnw/ni , \Urnw/nh , 
        \Uerr/nl , \Uerr/ni , \Uerr/nh , n1, n2, n6;
    assign \tc_wd[63]  = tc_wd[63];
    assign \tc_wd[62]  = tc_wd[62];
    assign \tc_wd[61]  = tc_wd[61];
    assign \tc_wd[60]  = tc_wd[60];
    assign \tc_wd[59]  = tc_wd[59];
    assign \tc_wd[58]  = tc_wd[58];
    assign \tc_wd[56]  = tc_wd[56];
    assign \tc_wd[55]  = tc_wd[55];
    assign \tc_wd[54]  = tc_wd[54];
    assign \tc_wd[53]  = tc_wd[53];
    assign \tc_wd[52]  = tc_wd[52];
    assign \tc_wd[51]  = tc_wd[51];
    assign \tc_wd[50]  = tc_wd[50];
    assign \tc_wd[49]  = tc_wd[49];
    assign \tc_wd[48]  = tc_wd[48];
    assign \tc_wd[47]  = tc_wd[47];
    assign \tc_wd[46]  = tc_wd[46];
    assign \tc_wd[45]  = tc_wd[45];
    assign \tc_wd[44]  = tc_wd[44];
    assign \tc_wd[43]  = tc_wd[43];
    assign \tc_wd[40]  = tc_wd[40];
    assign \tc_wd[39]  = tc_wd[39];
    assign \tc_wd[38]  = tc_wd[38];
    assign \tc_wd[36]  = tc_wd[36];
    assign \tc_wd[32]  = tc_wd[32];
    assign \tc_a[60]  = tc_a[60];
    assign \tc_a[58]  = tc_a[58];
    assign ts_i[2] = 1'b0;
    assign ts_i[1] = 1'b0;
    assign ts_i[0] = 1'b0;
    assign adr_i[28] = \tc_a[60] ;
    assign adr_i[26] = \tc_a[58] ;
    assign dat_i[31] = \tc_wd[63] ;
    assign dat_i[30] = \tc_wd[62] ;
    assign dat_i[29] = \tc_wd[61] ;
    assign dat_i[28] = \tc_wd[60] ;
    assign dat_i[27] = \tc_wd[59] ;
    assign dat_i[26] = \tc_wd[58] ;
    assign dat_i[24] = \tc_wd[56] ;
    assign dat_i[23] = \tc_wd[55] ;
    assign dat_i[22] = \tc_wd[54] ;
    assign dat_i[21] = \tc_wd[53] ;
    assign dat_i[20] = \tc_wd[52] ;
    assign dat_i[19] = \tc_wd[51] ;
    assign dat_i[18] = \tc_wd[50] ;
    assign dat_i[17] = \tc_wd[49] ;
    assign dat_i[16] = \tc_wd[48] ;
    assign dat_i[15] = \tc_wd[47] ;
    assign dat_i[14] = \tc_wd[46] ;
    assign dat_i[13] = \tc_wd[45] ;
    assign dat_i[12] = \tc_wd[44] ;
    assign dat_i[11] = \tc_wd[43] ;
    assign dat_i[8] = \tc_wd[40] ;
    assign dat_i[7] = \tc_wd[39] ;
    assign dat_i[6] = \tc_wd[38] ;
    assign dat_i[4] = \tc_wd[36] ;
    assign dat_i[0] = \tc_wd[32] ;
    assign prd_i = 1'b0;
    assign sel_i[3] = \sel_i[2] ;
    assign sel_i[2] = \sel_i[2] ;
    assign sel_i[0] = 1'b1;
    assign tc_ack = ack_in;
    assign ack_out = tr_ack;
    sr2dr_word_7 Urd ( .i(dat_o), .req(n2), .h(tr_rd[63:32]), .l(tr_rd[31:0])
         );
    inv_1 U3 ( .x(n334), .a(tc_a[7]) );
    inv_1 U5 ( .x(n311), .a(tc_a[21]) );
    and2_1 U6 ( .x(n129), .a(n309), .b(n310) );
    inv_1 U7 ( .x(n309), .a(tc_a[6]) );
    inv_1 U9 ( .x(n315), .a(tc_itag[4]) );
    nand2_1 U10 ( .x(n348), .a(n349), .b(n350) );
    inv_1 U11 ( .x(n349), .a(tc_a[12]) );
    inv_1 U12 ( .x(n456), .a(n348) );
    inv_1 U13 ( .x(n336), .a(tc_a[30]) );
    inv_1 U14 ( .x(n457), .a(n345) );
    inv_1 U15 ( .x(n303), .a(tc_a[8]) );
    nand3_1 U16 ( .x(n505), .a(n193), .b(n476), .c(n479) );
    inv_1 U17 ( .x(n229), .a(tc_wd[5]) );
    inv_1 U18 ( .x(n226), .a(tc_wd[3]) );
    inv_1 U19 ( .x(n257), .a(tc_wd[16]) );
    inv_1 U20 ( .x(n263), .a(tc_wd[21]) );
    inv_1 U21 ( .x(n260), .a(tc_wd[19]) );
    nand2_1 U22 ( .x(n268), .a(n269), .b(n270) );
    inv_1 U23 ( .x(n269), .a(tc_wd[23]) );
    inv_1 U24 ( .x(n270), .a(\tc_wd[55] ) );
    nand2_1 U25 ( .x(n265), .a(n266), .b(n267) );
    inv_1 U26 ( .x(n266), .a(tc_wd[20]) );
    inv_1 U27 ( .x(n277), .a(tc_wd[27]) );
    inv_1 U28 ( .x(n252), .a(\tc_wd[47] ) );
    nand2_1 U29 ( .x(n248), .a(n249), .b(n250) );
    inv_1 U30 ( .x(n249), .a(tc_wd[12]) );
    nand2_1 U31 ( .x(n245), .a(n246), .b(n247) );
    inv_1 U32 ( .x(n246), .a(tc_wd[13]) );
    inv_1 U33 ( .x(n247), .a(\tc_wd[45] ) );
    nand2_1 U34 ( .x(n242), .a(n243), .b(n244) );
    inv_1 U35 ( .x(n243), .a(tc_wd[11]) );
    nand2_1 U36 ( .x(n222), .a(n223), .b(n224) );
    inv_1 U37 ( .x(n223), .a(tc_wd[0]) );
    inv_1 U38 ( .x(n220), .a(tc_wd[1]) );
    nand2_1 U39 ( .x(n234), .a(n235), .b(n236) );
    inv_1 U40 ( .x(n235), .a(tc_wd[7]) );
    nand2_1 U41 ( .x(n231), .a(n232), .b(n233) );
    inv_1 U42 ( .x(n232), .a(tc_wd[4]) );
    nand2_1 U43 ( .x(n205), .a(n206), .b(n207) );
    inv_1 U44 ( .x(n206), .a(tc_wd[18]) );
    inv_1 U45 ( .x(n203), .a(tc_wd[10]) );
    nand2_1 U46 ( .x(n199), .a(n200), .b(n201) );
    inv_1 U47 ( .x(n200), .a(tc_wd[6]) );
    inv_1 U48 ( .x(n197), .a(tc_wd[2]) );
    inv_1 U49 ( .x(n218), .a(\tc_wd[46] ) );
    nand2_1 U50 ( .x(n214), .a(n215), .b(n216) );
    inv_1 U51 ( .x(n215), .a(tc_wd[30]) );
    nand2_1 U52 ( .x(n211), .a(n212), .b(n213) );
    inv_1 U53 ( .x(n213), .a(\tc_wd[58] ) );
    nand2_1 U54 ( .x(n208), .a(n209), .b(n210) );
    inv_1 U55 ( .x(n209), .a(tc_wd[22]) );
    inv_1 U56 ( .x(n374), .a(tc_rnw[0]) );
    inv_1 U57 ( .x(n375), .a(tc_rnw[1]) );
    inv_1 U58 ( .x(n368), .a(tc_a[18]) );
    inv_1 U59 ( .x(n244), .a(\tc_wd[43] ) );
    inv_1 U60 ( .x(n251), .a(tc_wd[15]) );
    inv_1 U61 ( .x(n250), .a(\tc_wd[44] ) );
    inv_1 U62 ( .x(n280), .a(tc_wd[29]) );
    inv_1 U63 ( .x(n267), .a(\tc_wd[52] ) );
    inv_1 U64 ( .x(n274), .a(tc_wd[24]) );
    inv_1 U65 ( .x(n271), .a(tc_wd[25]) );
    inv_1 U66 ( .x(n212), .a(tc_wd[26]) );
    inv_1 U67 ( .x(n210), .a(\tc_wd[54] ) );
    inv_1 U68 ( .x(n216), .a(\tc_wd[62] ) );
    inv_1 U69 ( .x(n201), .a(\tc_wd[38] ) );
    inv_1 U70 ( .x(n427), .a(n196) );
    inv_1 U71 ( .x(n207), .a(\tc_wd[50] ) );
    inv_1 U72 ( .x(n424), .a(n202) );
    inv_1 U73 ( .x(n236), .a(\tc_wd[39] ) );
    inv_1 U74 ( .x(n233), .a(\tc_wd[36] ) );
    inv_1 U75 ( .x(n240), .a(tc_wd[8]) );
    inv_1 U76 ( .x(n237), .a(tc_wd[9]) );
    inv_1 U77 ( .x(n224), .a(\tc_wd[32] ) );
    inv_1 U78 ( .x(n413), .a(n219) );
    nand2_1 U79 ( .x(n421), .a(n418), .b(n416) );
    nand2_1 U80 ( .x(n428), .a(n425), .b(n422) );
    nand2_1 U81 ( .x(n414), .a(n411), .b(n408) );
    inv_1 U82 ( .x(n238), .a(tc_wd[41]) );
    inv_1 U83 ( .x(n272), .a(tc_wd[57]) );
    inv_1 U84 ( .x(n350), .a(tc_a[44]) );
    inv_1 U85 ( .x(n351), .a(tc_a[43]) );
    inv_1 U86 ( .x(n366), .a(tc_a[41]) );
    inv_1 U87 ( .x(n335), .a(tc_a[39]) );
    inv_1 U88 ( .x(n310), .a(tc_a[38]) );
    inv_1 U89 ( .x(n355), .a(tc_a[52]) );
    and3_1 U90 ( .x(tc_ok), .a(n531), .b(n532), .c(respond) );
    and2_1 U91 ( .x(tc_slow), .a(respond), .b(acc_o) );
    inv_1 U94 ( .x(n313), .a(tc_itag[5]) );
    and2_1 U95 ( .x(n121), .a(n334), .b(n335) );
    and2_1 U96 ( .x(n122), .a(n359), .b(n360) );
    and2_1 U97 ( .x(n123), .a(n336), .b(n337) );
    and2_1 U98 ( .x(n124), .a(n237), .b(n238) );
    and2_1 U99 ( .x(n125), .a(n251), .b(n252) );
    and2_1 U100 ( .x(n126), .a(n271), .b(n272) );
    and2_1 U101 ( .x(n127), .a(n217), .b(n218) );
    and2_1 U102 ( .x(n128), .a(n311), .b(n312) );
    nor2_1 U103 ( .x(n130), .a(n1), .b(tc_size[2]) );
    nand2i_1 U105 ( .x(n284), .a(tc_wd[31]), .b(n285) );
    oa22_1 U106 ( .x(n449), .a(tc_a[27]), .b(tc_a[59]), .c(tc_a[54]), .d(tc_a
        [22]) );
    inv_1 U107 ( .x(n359), .a(tc_a[27]) );
    inv_1 U108 ( .x(n360), .a(tc_a[59]) );
    nand2i_1 U109 ( .x(n282), .a(tc_wd[28]), .b(n283) );
    nor2_1 U110 ( .x(n479), .a(tc_itag[0]), .b(tc_itag[5]) );
    nand4_1 U112 ( .x(n380), .a(n279), .b(n276), .c(n284), .d(n282) );
    aoi21_1 U113 ( .x(n425), .a(n200), .b(n201), .c(n427) );
    oa22_1 U114 ( .x(n397), .a(tc_wd[13]), .b(\tc_wd[45] ), .c(tc_wd[11]), .d(
        \tc_wd[43] ) );
    nor2_1 U115 ( .x(n454), .a(tc_a[20]), .b(tc_a[52]) );
    aoi21_1 U116 ( .x(n422), .a(n206), .b(n207), .c(n424) );
    oa22_1 U117 ( .x(n418), .a(tc_wd[26]), .b(\tc_wd[58] ), .c(tc_wd[22]), .d(
        \tc_wd[54] ) );
    oa22_1 U118 ( .x(n416), .a(tc_wd[14]), .b(\tc_wd[46] ), .c(tc_wd[30]), .d(
        \tc_wd[62] ) );
    inv_1 U119 ( .x(n217), .a(tc_wd[14]) );
    aoi22_1 U120 ( .x(n463), .a(n336), .b(n337), .c(n334), .d(n335) );
    nor2_1 U121 ( .x(n453), .a(tc_a[11]), .b(tc_a[43]) );
    oa22_1 U122 ( .x(n395), .a(tc_wd[15]), .b(\tc_wd[47] ), .c(tc_wd[12]), .d(
        \tc_wd[44] ) );
    oa22_1 U123 ( .x(n404), .a(tc_wd[7]), .b(\tc_wd[39] ), .c(tc_wd[4]), .d(
        \tc_wd[36] ) );
    oa22_1 U124 ( .x(n383), .a(tc_wd[23]), .b(\tc_wd[55] ), .c(tc_wd[20]), .d(
        \tc_wd[52] ) );
    aoi21_1 U125 ( .x(n411), .a(n223), .b(n224), .c(n413) );
    nor2_1 U126 ( .x(n443), .a(tc_a[49]), .b(tc_a[17]) );
    aoi22_1 U127 ( .x(n477), .a(n311), .b(n312), .c(n309), .d(n310) );
    oa21_1 U128 ( .x(n455), .a(tc_a[12]), .b(tc_a[44]), .c(n345) );
    inv_1 U129 ( .x(dat_i[5]), .a(n230) );
    inv_1 U130 ( .x(dat_i[9]), .a(n238) );
    inv_1 U131 ( .x(dat_i[25]), .a(n272) );
    buf_1 U132 ( .x(\sel_i[2] ), .a(n1) );
    buf_1 U133 ( .x(adr_i[16]), .a(tc_a[48]) );
    nor2_1 U134 ( .x(n135), .a(tc_a[14]), .b(tc_a[46]) );
    inv_1 U135 ( .x(n305), .a(tc_a[46]) );
    inv_1 U136 ( .x(n487), .a(n302) );
    nand2i_1 U137 ( .x(n445), .a(n446), .b(n442) );
    nor2_1 U138 ( .x(n136), .a(tc_a[29]), .b(tc_a[61]) );
    inv_1 U139 ( .x(n320), .a(tc_a[61]) );
    nand2_1 U140 ( .x(n400), .a(n397), .b(n395) );
    inv_1 U141 ( .x(n137), .a(n340) );
    inv_1 U142 ( .x(dat_i[2]), .a(n198) );
    nand2_1 U143 ( .x(n386), .a(n383), .b(n381) );
    nand3i_1 U144 ( .x(n478), .a(n479), .b(n477), .c(n475) );
    nand2_1 U145 ( .x(n407), .a(n404), .b(n402) );
    inv_1 U146 ( .x(dat_i[10]), .a(n204) );
    inv_1 U147 ( .x(dat_i[1]), .a(n221) );
    nor2_1 U148 ( .x(n141), .a(tc_a[3]), .b(tc_a[35]) );
    inv_1 U149 ( .x(n321), .a(tc_a[35]) );
    nor2_1 U151 ( .x(n483), .a(n484), .b(n485) );
    nor2_1 U152 ( .x(n480), .a(n474), .b(n478) );
    inv_1 U153 ( .x(dat_i[3]), .a(n227) );
    nor2_1 U154 ( .x(n188), .a(n517), .b(n525) );
    nand2_1 U155 ( .x(n180), .a(n401), .b(n387) );
    nor2_1 U156 ( .x(n401), .a(n394), .b(n400) );
    nor2_1 U157 ( .x(n387), .a(n380), .b(n386) );
    nor2_1 U158 ( .x(n481), .a(n482), .b(n135) );
    nor2_1 U159 ( .x(n491), .a(n195), .b(n492) );
    nor2_1 U160 ( .x(n195), .a(tc_size[1]), .b(n1) );
    inv_1 U161 ( .x(adr_i[18]), .a(n369) );
    nand2_1 U162 ( .x(n181), .a(n429), .b(n415) );
    nor2_1 U163 ( .x(n429), .a(n421), .b(n428) );
    nor2_1 U164 ( .x(n415), .a(n407), .b(n414) );
    inv_1 U165 ( .x(adr_i[0]), .a(n324) );
    inv_1 U166 ( .x(n324), .a(tc_a[32]) );
    inv_1 U167 ( .x(sel_i[1]), .a(n130) );
    inv_1 U168 ( .x(st_i[2]), .a(n343) );
    inv_1 U169 ( .x(adr_i[9]), .a(n366) );
    inv_1 U170 ( .x(adr_i[24]), .a(n363) );
    inv_1 U171 ( .x(adr_i[19]), .a(n319) );
    inv_1 U172 ( .x(n319), .a(tc_a[51]) );
    inv_1 U173 ( .x(n369), .a(tc_a[50]) );
    inv_1 U174 ( .x(st_i[3]), .a(n344) );
    inv_1 U175 ( .x(adr_i[13]), .a(n354) );
    inv_1 U176 ( .x(adr_i[12]), .a(n350) );
    inv_1 U177 ( .x(adr_i[8]), .a(n304) );
    inv_1 U178 ( .x(n304), .a(tc_a[40]) );
    inv_1 U179 ( .x(adr_i[2]), .a(n330) );
    buf_1 U180 ( .x(adr_i[17]), .a(tc_a[49]) );
    nand2_1 U181 ( .x(n497), .a(n496), .b(n130) );
    inv_1 U182 ( .x(adr_i[10]), .a(n291) );
    and2_1 U183 ( .x(n438), .a(n373), .b(n367) );
    inv_1 U184 ( .x(n439), .a(n373) );
    inv_1 U185 ( .x(n440), .a(n367) );
    inv_1 U186 ( .x(adr_i[20]), .a(n355) );
    inv_1 U187 ( .x(adr_i[27]), .a(n360) );
    inv_1 U188 ( .x(adr_i[4]), .a(n333) );
    inv_1 U189 ( .x(adr_i[25]), .a(n308) );
    inv_1 U190 ( .x(adr_i[30]), .a(n337) );
    inv_1 U191 ( .x(adr_i[31]), .a(n297) );
    inv_1 U192 ( .x(n297), .a(tc_a[63]) );
    inv_1 U193 ( .x(adr_i[15]), .a(n347) );
    inv_1 U194 ( .x(adr_i[11]), .a(n351) );
    inv_1 U195 ( .x(adr_i[1]), .a(n301) );
    inv_1 U196 ( .x(n301), .a(tc_a[33]) );
    nand2_1 U197 ( .x(n503), .a(n499), .b(n502) );
    nor2_1 U198 ( .x(n499), .a(n497), .b(n498) );
    inv_1 U199 ( .x(adr_i[21]), .a(n312) );
    inv_1 U200 ( .x(n312), .a(tc_a[53]) );
    inv_1 U201 ( .x(seq_i), .a(n288) );
    inv_1 U202 ( .x(adr_i[5]), .a(n327) );
    inv_1 U203 ( .x(st_i[4]), .a(n316) );
    inv_1 U204 ( .x(n316), .a(tc_itag[9]) );
    inv_1 U205 ( .x(st_i[1]), .a(n298) );
    inv_1 U206 ( .x(adr_i[23]), .a(n294) );
    inv_1 U207 ( .x(adr_i[22]), .a(n358) );
    nand2_1 U208 ( .x(complb0), .a(n188), .b(n189) );
    nor2_1 U209 ( .x(n189), .a(n503), .b(n510) );
    inv_1 U210 ( .x(adr_i[29]), .a(n320) );
    inv_1 U211 ( .x(adr_i[7]), .a(n335) );
    inv_1 U212 ( .x(adr_i[14]), .a(n305) );
    inv_1 U213 ( .x(adr_i[6]), .a(n310) );
    inv_1 U214 ( .x(st_i[0]), .a(n313) );
    inv_1 U215 ( .x(adr_i[3]), .a(n321) );
    nand3_1 U218 ( .x(n507), .a(n192), .b(n136), .c(n473) );
    nand2_1 U219 ( .x(n508), .a(n471), .b(n141) );
    nor2_1 U220 ( .x(n488), .a(n489), .b(n490) );
    nand4_1 U222 ( .x(complw0), .a(n182), .b(n183), .c(n184), .d(n185) );
    nor2_1 U223 ( .x(n192), .a(\tc_a[58] ), .b(tc_a[26]) );
    nor2_1 U224 ( .x(n193), .a(tc_a[48]), .b(tc_a[16]) );
    nand2_1 U225 ( .x(n364), .a(n365), .b(n366) );
    nand2_1 U226 ( .x(n394), .a(n391), .b(n388) );
    nand4_1 U227 ( .x(n430), .a(n423), .b(n424), .c(n426), .d(n427) );
    nand4_1 U228 ( .x(n431), .a(n127), .b(n417), .c(n419), .d(n420) );
    nor2_1 U229 ( .x(n185), .a(n430), .b(n431) );
    nand4_1 U230 ( .x(n432), .a(n409), .b(n410), .c(n412), .d(n413) );
    nand4_1 U231 ( .x(n433), .a(n403), .b(n124), .c(n405), .d(n406) );
    nor2_1 U232 ( .x(n184), .a(n432), .b(n433) );
    nand4_1 U233 ( .x(n434), .a(n125), .b(n396), .c(n398), .d(n399) );
    nand4_1 U234 ( .x(n435), .a(n389), .b(n390), .c(n392), .d(n393) );
    nor2_1 U235 ( .x(n183), .a(n434), .b(n435) );
    nand4_1 U236 ( .x(n436), .a(n382), .b(n126), .c(n384), .d(n385) );
    nand4_1 U237 ( .x(n437), .a(n376), .b(n377), .c(n378), .d(n379) );
    nor2_1 U238 ( .x(n182), .a(n436), .b(n437) );
    nand2_1 U239 ( .x(n441), .a(n438), .b(n370) );
    nor2_1 U240 ( .x(n442), .a(n443), .b(n444) );
    nor3_1 U241 ( .x(n470), .a(n471), .b(n136), .c(n141) );
    nor3_1 U242 ( .x(n472), .a(n473), .b(n192), .c(n193) );
    nand2_1 U243 ( .x(n474), .a(n472), .b(n470) );
    nor2_1 U244 ( .x(n475), .a(n476), .b(n194) );
    nand3i_1 U245 ( .x(n486), .a(n487), .b(n481), .c(n483) );
    nand3i_1 U246 ( .x(n493), .a(n494), .b(n488), .c(n491) );
    nor2_1 U247 ( .x(n495), .a(n493), .b(n486) );
    nand2_1 U248 ( .x(n191), .a(n495), .b(n480) );
    nand3_1 U249 ( .x(n498), .a(n489), .b(n492), .c(n490) );
    nand3_1 U250 ( .x(n500), .a(n485), .b(n494), .c(n484) );
    nand2_1 U251 ( .x(n501), .a(n135), .b(n487) );
    nor2_1 U252 ( .x(n502), .a(n500), .b(n501) );
    nand3_1 U253 ( .x(n504), .a(n128), .b(n482), .c(n129) );
    nor2_1 U254 ( .x(n506), .a(n504), .b(n505) );
    nor2_1 U255 ( .x(n509), .a(n507), .b(n508) );
    nand2_1 U256 ( .x(n510), .a(n509), .b(n506) );
    nand3_1 U257 ( .x(n511), .a(n465), .b(n466), .c(n468) );
    nand3_1 U258 ( .x(n512), .a(n123), .b(n121), .c(n460) );
    nor2_1 U259 ( .x(n513), .a(n511), .b(n512) );
    nand3_1 U260 ( .x(n514), .a(n462), .b(n459), .c(n457) );
    nand2_1 U261 ( .x(n515), .a(n453), .b(n456) );
    nor2_1 U262 ( .x(n516), .a(n514), .b(n515) );
    nand2_1 U263 ( .x(n517), .a(n516), .b(n513) );
    nand2_1 U264 ( .x(n518), .a(n454), .b(n452) );
    nor2i_1 U265 ( .x(n519), .a(n450), .b(n518) );
    nand2_1 U266 ( .x(n520), .a(n444), .b(n122) );
    nor2i_1 U267 ( .x(n522), .a(n446), .b(n521) );
    nand2_1 U268 ( .x(n523), .a(n439), .b(n524) );
    inv_1 U270 ( .x(n365), .a(tc_a[9]) );
    inv_1 U271 ( .x(n371), .a(\tc_a[60] ) );
    inv_1 U272 ( .x(n446), .a(n364) );
    nor2_1 U273 ( .x(complb1), .a(n190), .b(n191) );
    nor2_1 U274 ( .x(complw1), .a(n180), .b(n181) );
    nand3i_1 U276 ( .x(n190), .a(n441), .b(n447), .c(n469) );
    and4_1 U277 ( .x(n5), .a(n3), .b(n4), .c(n519), .d(n522) );
    inv_1 U216 ( .x(n3), .a(n520) );
    inv_1 U217 ( .x(n4), .a(n523) );
    inv_1 U428 ( .x(n525), .a(n5) );
    nor2_1 U278 ( .x(n447), .a(n448), .b(n445) );
    nor2_1 U279 ( .x(n469), .a(n467), .b(n461) );
    nand2_1 U280 ( .x(n370), .a(n371), .b(n372) );
    nand3i_1 U281 ( .x(n448), .a(n454), .b(n449), .c(n451) );
    nand3i_1 U282 ( .x(n461), .a(n462), .b(n455), .c(n458) );
    nand3i_1 U283 ( .x(n467), .a(n468), .b(n463), .c(n464) );
    inv_1 U284 ( .x(n382), .a(n273) );
    inv_1 U285 ( .x(n384), .a(n268) );
    inv_1 U286 ( .x(n385), .a(n265) );
    inv_1 U287 ( .x(n376), .a(n284) );
    inv_1 U288 ( .x(n377), .a(n282) );
    inv_1 U289 ( .x(n378), .a(n279) );
    inv_1 U290 ( .x(n379), .a(n276) );
    inv_1 U291 ( .x(n396), .a(n248) );
    inv_1 U292 ( .x(n398), .a(n245) );
    inv_1 U293 ( .x(n399), .a(n242) );
    inv_1 U294 ( .x(n389), .a(n262) );
    inv_1 U295 ( .x(n390), .a(n259) );
    inv_1 U296 ( .x(n392), .a(n256) );
    inv_1 U297 ( .x(n393), .a(n253) );
    inv_1 U298 ( .x(n409), .a(n228) );
    inv_1 U299 ( .x(n410), .a(n225) );
    inv_1 U300 ( .x(n412), .a(n222) );
    inv_1 U301 ( .x(n403), .a(n239) );
    inv_1 U302 ( .x(n405), .a(n234) );
    inv_1 U303 ( .x(n406), .a(n231) );
    inv_1 U304 ( .x(n423), .a(n205) );
    inv_1 U305 ( .x(n426), .a(n199) );
    inv_1 U306 ( .x(n417), .a(n214) );
    inv_1 U307 ( .x(n419), .a(n211) );
    inv_1 U308 ( .x(n420), .a(n208) );
    inv_1 U309 ( .x(n444), .a(n361) );
    inv_1 U310 ( .x(n524), .a(n370) );
    inv_1 U311 ( .x(n450), .a(n356) );
    nand2_1 U312 ( .x(n521), .a(n443), .b(n440) );
    inv_1 U313 ( .x(n372), .a(tc_a[28]) );
    nor2_1 U314 ( .x(n451), .a(n452), .b(n453) );
    nor2_1 U315 ( .x(n458), .a(n459), .b(n460) );
    inv_1 U316 ( .x(n468), .a(n331) );
    nor2_1 U317 ( .x(n464), .a(n465), .b(n466) );
    inv_1 U318 ( .x(n494), .a(n295) );
    nand2_1 U319 ( .x(n273), .a(n274), .b(n275) );
    nand2_1 U320 ( .x(n279), .a(n280), .b(n281) );
    nand2_1 U321 ( .x(n276), .a(n277), .b(n278) );
    nand2_1 U322 ( .x(n262), .a(n263), .b(n264) );
    nand2_1 U323 ( .x(n259), .a(n260), .b(n261) );
    nand2_1 U324 ( .x(n256), .a(n257), .b(n258) );
    nand2_1 U325 ( .x(n253), .a(n254), .b(n255) );
    nand2_1 U326 ( .x(n228), .a(n229), .b(n230) );
    nand2_1 U327 ( .x(n225), .a(n226), .b(n227) );
    nand2_1 U328 ( .x(n219), .a(n220), .b(n221) );
    nand2_1 U329 ( .x(n239), .a(n240), .b(n241) );
    nand2_1 U330 ( .x(n202), .a(n203), .b(n204) );
    nand2_1 U331 ( .x(n196), .a(n197), .b(n198) );
    nor2_1 U332 ( .x(n391), .a(n392), .b(n393) );
    nor2_1 U333 ( .x(n388), .a(n389), .b(n390) );
    nor2_1 U334 ( .x(n381), .a(n382), .b(n126) );
    nor2_1 U335 ( .x(n402), .a(n403), .b(n124) );
    nor2_1 U336 ( .x(n408), .a(n409), .b(n410) );
    inv_1 U337 ( .x(n459), .a(n341) );
    inv_1 U338 ( .x(n465), .a(n328) );
    inv_1 U339 ( .x(n466), .a(n325) );
    inv_1 U340 ( .x(n460), .a(n338) );
    nand2_1 U341 ( .x(n361), .a(n362), .b(n363) );
    nand2_1 U342 ( .x(n373), .a(n374), .b(n375) );
    nand2_1 U343 ( .x(n356), .a(n358), .b(n357) );
    inv_1 U344 ( .x(n452), .a(n352) );
    inv_1 U345 ( .x(n484), .a(n299) );
    inv_1 U346 ( .x(n489), .a(n289) );
    inv_1 U347 ( .x(n492), .a(n286) );
    inv_1 U348 ( .x(n490), .a(n292) );
    inv_1 U349 ( .x(n473), .a(n317) );
    inv_1 U350 ( .x(n471), .a(n322) );
    inv_1 U351 ( .x(n482), .a(n306) );
    inv_1 U352 ( .x(n476), .a(n314) );
    nand2_1 U353 ( .x(n367), .a(n368), .b(n369) );
    nand2_1 U354 ( .x(n331), .a(n332), .b(n333) );
    nand2_1 U355 ( .x(n302), .a(n303), .b(n304) );
    nand2_1 U356 ( .x(n295), .a(n296), .b(n297) );
    inv_1 U357 ( .x(n275), .a(\tc_wd[56] ) );
    inv_1 U358 ( .x(n285), .a(\tc_wd[63] ) );
    inv_1 U359 ( .x(n283), .a(\tc_wd[60] ) );
    inv_1 U360 ( .x(n281), .a(\tc_wd[61] ) );
    inv_1 U361 ( .x(n278), .a(\tc_wd[59] ) );
    inv_1 U362 ( .x(n264), .a(\tc_wd[53] ) );
    inv_1 U363 ( .x(n261), .a(\tc_wd[51] ) );
    inv_1 U364 ( .x(n258), .a(\tc_wd[48] ) );
    inv_1 U365 ( .x(n254), .a(tc_wd[17]) );
    inv_1 U366 ( .x(n255), .a(\tc_wd[49] ) );
    inv_1 U367 ( .x(n230), .a(tc_wd[37]) );
    inv_1 U368 ( .x(n227), .a(tc_wd[35]) );
    inv_1 U369 ( .x(n221), .a(tc_wd[33]) );
    inv_1 U370 ( .x(n241), .a(\tc_wd[40] ) );
    inv_1 U371 ( .x(n204), .a(tc_wd[42]) );
    inv_1 U372 ( .x(n198), .a(tc_wd[34]) );
    nand2_1 U373 ( .x(n341), .a(n342), .b(n343) );
    nand2_1 U374 ( .x(n345), .a(n347), .b(n346) );
    nand2_1 U375 ( .x(n328), .a(n329), .b(n330) );
    nand2_1 U376 ( .x(n325), .a(n326), .b(n327) );
    nand2_1 U377 ( .x(n338), .a(n340), .b(n339) );
    inv_1 U378 ( .x(n362), .a(tc_a[24]) );
    inv_1 U379 ( .x(n363), .a(tc_a[56]) );
    inv_1 U380 ( .x(n357), .a(tc_a[22]) );
    inv_1 U381 ( .x(n358), .a(tc_a[54]) );
    nand2_1 U382 ( .x(n352), .a(n353), .b(n354) );
    nand2_1 U383 ( .x(n299), .a(n300), .b(n301) );
    nand2_1 U384 ( .x(n289), .a(n290), .b(n291) );
    nand2_1 U385 ( .x(n286), .a(n287), .b(n288) );
    nand2_1 U386 ( .x(n292), .a(n293), .b(n294) );
    nand2_1 U387 ( .x(n317), .a(n318), .b(n319) );
    nand2_1 U388 ( .x(n322), .a(n323), .b(n324) );
    nand2_1 U389 ( .x(n306), .a(n307), .b(n308) );
    nand2_1 U390 ( .x(n314), .a(n315), .b(n316) );
    inv_1 U391 ( .x(n332), .a(tc_a[4]) );
    inv_1 U392 ( .x(n333), .a(tc_a[36]) );
    inv_1 U393 ( .x(n296), .a(tc_a[31]) );
    inv_1 U394 ( .x(n342), .a(tc_itag[2]) );
    inv_1 U395 ( .x(n343), .a(tc_itag[7]) );
    inv_1 U396 ( .x(n346), .a(tc_a[15]) );
    inv_1 U397 ( .x(n347), .a(tc_a[47]) );
    inv_1 U398 ( .x(n329), .a(tc_a[2]) );
    inv_1 U399 ( .x(n330), .a(tc_a[34]) );
    inv_1 U400 ( .x(n326), .a(tc_a[5]) );
    inv_1 U401 ( .x(n327), .a(tc_a[37]) );
    inv_1 U402 ( .x(n337), .a(tc_a[62]) );
    inv_1 U403 ( .x(n339), .a(tc_lock[0]) );
    inv_1 U404 ( .x(n340), .a(tc_lock[1]) );
    inv_1 U405 ( .x(n353), .a(tc_a[13]) );
    inv_1 U406 ( .x(n354), .a(tc_a[45]) );
    inv_1 U407 ( .x(n300), .a(tc_a[1]) );
    inv_1 U408 ( .x(n290), .a(tc_a[10]) );
    inv_1 U409 ( .x(n291), .a(tc_a[42]) );
    inv_1 U410 ( .x(n287), .a(tc_seq[0]) );
    inv_1 U411 ( .x(n288), .a(tc_seq[1]) );
    inv_1 U412 ( .x(n293), .a(tc_a[23]) );
    inv_1 U413 ( .x(n294), .a(tc_a[55]) );
    inv_1 U414 ( .x(n318), .a(tc_a[19]) );
    inv_1 U415 ( .x(n323), .a(tc_a[0]) );
    inv_1 U416 ( .x(n307), .a(tc_a[25]) );
    inv_1 U417 ( .x(n308), .a(tc_a[57]) );
    buf_1 U418 ( .x(we_i), .a(tc_rnw[0]) );
    matched_delay_cp2slave_resp_imem U419 ( .x(req_out_delayed), .a(req_out)
         );
    and4_1 U420 ( .x(_25_net_), .a(sel_o[0]), .b(sel_o[1]), .c(n529), .d(n530)
         );
    inv_1 U421 ( .x(_24_net_), .a(we_i) );
    and2_1 U422 ( .x(tc_defer), .a(rty_o), .b(respond) );
    and4_1 U423 ( .x(_26_net_), .a(sel_o[0]), .b(sel_o[1]), .c(sel_o[3]), .d(
        sel_o[2]) );
    inv_1 U424 ( .x(n532), .a(acc_o) );
    inv_1 U425 ( .x(n531), .a(rty_o) );
    inv_1 U426 ( .x(n529), .a(sel_o[2]) );
    inv_1 U427 ( .x(n530), .a(sel_o[3]) );
    buf_1 U150 ( .x(n142), .a(req_in_i) );
    matched_delay_cp2slave_comimem matchDelCom ( .x(req_in), .a(req_in_i) );
    nand2_1 U275 ( .x(req_in_i), .a(n186), .b(n187) );
    inv_1 U221 ( .x(n186), .a(all_w) );
    inv_1 U269 ( .x(n187), .a(all_r) );
    dffp_1 mult_i_reg ( .q(mult_i), .d(n137), .ck(n142) );
    ao222_1 \cg_respond/__tmp99/U1  ( .x(respond), .a(req_out), .b(tc_ack), 
        .c(req_out), .d(respond), .e(tc_ack), .f(respond) );
    oa21_1 \cg_all_r/__tmp99/U1  ( .x(all_r), .a(tc_rnw[1]), .b(all_r), .c(
        comp_basic) );
    ao31_1 \cg_all_w/__tmp99/aoi  ( .x(\cg_all_w/__tmp99/loop ), .a(comp_basic
        ), .b(comp_wd), .c(we_i), .d(all_w) );
    oa21_1 \cg_all_w/__tmp99/outGate  ( .x(all_w), .a(comp_basic), .b(comp_wd), 
        .c(\cg_all_w/__tmp99/loop ) );
    ao222_1 \cg_wd/__tmp99/U1  ( .x(comp_wd), .a(complw0), .b(complw1), .c(
        complw0), .d(comp_wd), .e(complw1), .f(comp_wd) );
    ao222_1 \cg_basic/__tmp99/U1  ( .x(comp_basic), .a(complb0), .b(complb1), 
        .c(complb0), .d(comp_basic), .e(complb1), .f(comp_basic) );
    inv_1 \Usze1/Uii  ( .x(\Usze1/ni ), .a(_26_net_) );
    inv_1 \Usze1/Uih  ( .x(\Usze1/nh ), .a(tr_size[3]) );
    inv_1 \Usze1/Uil  ( .x(\Usze1/nl ), .a(tr_size[1]) );
    ao23_1 \Usze1/Ucl/U1/U1  ( .x(tr_size[1]), .a(n6), .b(tr_size[1]), .c(n2), 
        .d(\Usze1/ni ), .e(\Usze1/nh ) );
    ao23_1 \Usze1/Uch/U1/U1  ( .x(tr_size[3]), .a(n2), .b(tr_size[3]), .c(n2), 
        .d(_26_net_), .e(\Usze1/nl ) );
    inv_1 \Usze0/Uii  ( .x(\Usze0/ni ), .a(_25_net_) );
    inv_1 \Usze0/Uih  ( .x(\Usze0/nh ), .a(tr_size[2]) );
    inv_1 \Usze0/Uil  ( .x(\Usze0/nl ), .a(tr_size[0]) );
    ao23_1 \Usze0/Ucl/U1/U1  ( .x(tr_size[0]), .a(n6), .b(tr_size[0]), .c(n2), 
        .d(\Usze0/ni ), .e(\Usze0/nh ) );
    ao23_1 \Usze0/Uch/U1/U1  ( .x(tr_size[2]), .a(n6), .b(tr_size[2]), .c(n2), 
        .d(_25_net_), .e(\Usze0/nl ) );
    inv_1 \Urnw/Uii  ( .x(\Urnw/ni ), .a(_24_net_) );
    inv_1 \Urnw/Uih  ( .x(\Urnw/nh ), .a(tr_rnw[1]) );
    inv_1 \Urnw/Uil  ( .x(\Urnw/nl ), .a(tr_rnw[0]) );
    ao23_1 \Urnw/Ucl/U1/U1  ( .x(tr_rnw[0]), .a(n2), .b(tr_rnw[0]), .c(n2), 
        .d(\Urnw/ni ), .e(\Urnw/nh ) );
    ao23_1 \Urnw/Uch/U1/U1  ( .x(tr_rnw[1]), .a(n2), .b(tr_rnw[1]), .c(n2), 
        .d(_24_net_), .e(\Urnw/nl ) );
    inv_1 \Uerr/Uii  ( .x(\Uerr/ni ), .a(err_o) );
    inv_1 \Uerr/Uih  ( .x(\Uerr/nh ), .a(tr_err[1]) );
    inv_1 \Uerr/Uil  ( .x(\Uerr/nl ), .a(tr_err[0]) );
    ao23_1 \Uerr/Ucl/U1/U1  ( .x(tr_err[0]), .a(n2), .b(tr_err[0]), .c(n2), 
        .d(\Uerr/ni ), .e(\Uerr/nh ) );
    ao23_1 \Uerr/Uch/U1/U1  ( .x(tr_err[1]), .a(n2), .b(tr_err[1]), .c(n2), 
        .d(err_o), .e(\Uerr/nl ) );
    inv_0 U1 ( .x(n344), .a(tc_itag[8]) );
    nor2_0 U2 ( .x(n462), .a(tc_itag[3]), .b(tc_itag[8]) );
    inv_0 U4 ( .x(n298), .a(tc_itag[6]) );
    nor2_0 U8 ( .x(n485), .a(tc_itag[1]), .b(tc_itag[6]) );
    nor2_0 U92 ( .x(n496), .a(tc_size[0]), .b(tc_size[1]) );
    nor2_0 U93 ( .x(n194), .a(tc_size[0]), .b(tc_size[2]) );
    buf_1 U104 ( .x(n1), .a(tc_size[3]) );
    buf_16 U111 ( .x(n2), .a(req_out_delayed) );
    buf_16 U429 ( .x(n6), .a(req_out_delayed) );
endmodule


module slave_if_imem ( nReset, sc_req, sc_we, sc_mult, sc_seq, sc_prd, sc_ts, 
    sc_st, sc_sel, sc_adr, sc_dat, sc_ack, sr_req, sr_err, sr_rty, sr_acc, 
    sr_mult, sr_ts, sr_rt, sr_sel, sr_dat, sr_ack, chaincommand, 
    nchaincommandack, chainresponse, nchainresponseack, e_dp, e_ip, e_tic, 
    r_dp, r_ip, r_tic );
output [2:0] sc_ts;
output [4:0] sc_st;
output [3:0] sc_sel;
output [31:0] sc_adr;
output [31:0] sc_dat;
input  [2:0] sr_ts;
input  [4:0] sr_rt;
input  [3:0] sr_sel;
input  [31:0] sr_dat;
input  [4:0] chaincommand;
output [4:0] chainresponse;
input  [2:0] e_dp;
input  [2:0] e_ip;
input  [2:0] e_tic;
input  [2:0] r_dp;
input  [2:0] r_ip;
input  [2:0] r_tic;
input  nReset, sc_ack, sr_req, sr_err, sr_rty, sr_acc, sr_mult, 
    nchainresponseack;
output sc_req, sc_we, sc_mult, sc_seq, sc_prd, sr_ack, nchaincommandack;
    wire \ct_a[63] , \ct_a[62] , \ct_a[61] , \ct_a[60] , \ct_a[59] , 
        \ct_a[58] , \ct_a[57] , \ct_a[56] , \ct_a[55] , \ct_a[54] , \ct_a[53] , 
        \ct_a[52] , \ct_a[51] , \ct_a[50] , \ct_a[49] , \ct_a[48] , \ct_a[47] , 
        \ct_a[46] , \ct_a[45] , \ct_a[44] , \ct_a[43] , \ct_a[42] , \ct_a[41] , 
        \ct_a[40] , \ct_a[39] , \ct_a[38] , \ct_a[37] , \ct_a[36] , \ct_a[35] , 
        \ct_a[34] , \ct_a[33] , \ct_a[32] , \ct_a[31] , \ct_a[30] , \ct_a[29] , 
        \ct_a[28] , \ct_a[27] , \ct_a[26] , \ct_a[25] , \ct_a[24] , \ct_a[23] , 
        \ct_a[22] , \ct_a[21] , \ct_a[20] , \ct_a[19] , \ct_a[18] , \ct_a[17] , 
        \ct_a[16] , \ct_a[15] , \ct_a[14] , \ct_a[13] , \ct_a[12] , \ct_a[11] , 
        \ct_a[10] , \ct_a[9] , \ct_a[8] , \ct_a[7] , \ct_a[6] , \ct_a[5] , 
        \ct_a[4] , \ct_a[3] , \ct_a[2] , \ct_a[1] , \ct_a[0] , \ct_wd[63] , 
        \ct_wd[62] , \ct_wd[61] , \ct_wd[60] , \ct_wd[59] , \ct_wd[58] , 
        \ct_wd[57] , \ct_wd[56] , \ct_wd[55] , \ct_wd[54] , \ct_wd[53] , 
        \ct_wd[52] , \ct_wd[51] , \ct_wd[50] , \ct_wd[49] , \ct_wd[48] , 
        \ct_wd[47] , \ct_wd[46] , \ct_wd[45] , \ct_wd[44] , \ct_wd[43] , 
        \ct_wd[42] , \ct_wd[41] , \ct_wd[40] , \ct_wd[39] , \ct_wd[38] , 
        \ct_wd[37] , \ct_wd[36] , \ct_wd[35] , \ct_wd[34] , \ct_wd[33] , 
        \ct_wd[32] , \ct_wd[31] , \ct_wd[30] , \ct_wd[29] , \ct_wd[28] , 
        \ct_wd[27] , \ct_wd[26] , \ct_wd[25] , \ct_wd[24] , \ct_wd[23] , 
        \ct_wd[22] , \ct_wd[21] , \ct_wd[20] , \ct_wd[19] , \ct_wd[18] , 
        \ct_wd[17] , \ct_wd[16] , \ct_wd[15] , \ct_wd[14] , \ct_wd[13] , 
        \ct_wd[12] , \ct_wd[11] , \ct_wd[10] , \ct_wd[9] , \ct_wd[8] , 
        \ct_wd[7] , \ct_wd[6] , \ct_wd[5] , \ct_wd[4] , \ct_wd[3] , \ct_wd[2] , 
        \ct_wd[1] , \ct_wd[0] , \ct_rnw[1] , \ct_rnw[0] , \ct_lock[1] , 
        \ct_lock[0] , \ct_seq[1] , \ct_seq[0] , \ct_size[3] , \ct_size[2] , 
        \ct_size[1] , \ct_size[0] , \ct_itag[9] , \ct_itag[8] , \ct_itag[7] , 
        \ct_itag[6] , \ct_itag[5] , \ct_itag[4] , \ct_itag[3] , \ct_itag[2] , 
        \ct_itag[1] , \ct_itag[0] , ct_ack, ct_ok, ct_defer, ct_slow, 
        \rt_rd[63] , \rt_rd[62] , \rt_rd[61] , \rt_rd[60] , \rt_rd[59] , 
        \rt_rd[58] , \rt_rd[57] , \rt_rd[56] , \rt_rd[55] , \rt_rd[54] , 
        \rt_rd[53] , \rt_rd[52] , \rt_rd[51] , \rt_rd[50] , \rt_rd[49] , 
        \rt_rd[48] , \rt_rd[47] , \rt_rd[46] , \rt_rd[45] , \rt_rd[44] , 
        \rt_rd[43] , \rt_rd[42] , \rt_rd[41] , \rt_rd[40] , \rt_rd[39] , 
        \rt_rd[38] , \rt_rd[37] , \rt_rd[36] , \rt_rd[35] , \rt_rd[34] , 
        \rt_rd[33] , \rt_rd[32] , \rt_rd[31] , \rt_rd[30] , \rt_rd[29] , 
        \rt_rd[28] , \rt_rd[27] , \rt_rd[26] , \rt_rd[25] , \rt_rd[24] , 
        \rt_rd[23] , \rt_rd[22] , \rt_rd[21] , \rt_rd[20] , \rt_rd[19] , 
        \rt_rd[18] , \rt_rd[17] , \rt_rd[16] , \rt_rd[15] , \rt_rd[14] , 
        \rt_rd[13] , \rt_rd[12] , \rt_rd[11] , \rt_rd[10] , \rt_rd[9] , 
        \rt_rd[8] , \rt_rd[7] , \rt_rd[6] , \rt_rd[5] , \rt_rd[4] , \rt_rd[3] , 
        \rt_rd[2] , \rt_rd[1] , \rt_rd[0] , \rt_err[1] , \rt_err[0] , rt_ack, 
        \tag_h[4] , \tag_h[3] , \tag_h[2] , \tag_h[1] , \tag_h[0] , \tag_l[4] , 
        \tag_l[3] , \tag_l[2] , \tag_l[1] , \tag_l[0] , \route[4] , \route[1] , 
        \route[0] , nroute_ack, routetx_req, routetx_ack, \eh[1] , \eh[0] , 
        \el[2] , \el[1] , \el[0] , \rh[2] , \rh[1] , \rl[2] , \rl[1] , \rl[0] , 
        reset;
    wire SYNOPSYS_UNCONNECTED_1 , SYNOPSYS_UNCONNECTED_2 , 
	SYNOPSYS_UNCONNECTED_3 , SYNOPSYS_UNCONNECTED_4 , SYNOPSYS_UNCONNECTED_5 ;
    assign sc_prd = 1'b0;
    assign sc_ts[2] = 1'b0;
    assign sc_ts[1] = 1'b0;
    assign sc_ts[0] = 1'b0;
    assign sc_sel[0] = 1'b1;
    target_imem tg ( .addr({\ct_a[63] , \ct_a[62] , \ct_a[61] , \ct_a[60] , 
        \ct_a[59] , \ct_a[58] , \ct_a[57] , \ct_a[56] , \ct_a[55] , \ct_a[54] , 
        \ct_a[53] , \ct_a[52] , \ct_a[51] , \ct_a[50] , \ct_a[49] , \ct_a[48] , 
        \ct_a[47] , \ct_a[46] , \ct_a[45] , \ct_a[44] , \ct_a[43] , \ct_a[42] , 
        \ct_a[41] , \ct_a[40] , \ct_a[39] , \ct_a[38] , \ct_a[37] , \ct_a[36] , 
        \ct_a[35] , \ct_a[34] , \ct_a[33] , \ct_a[32] , \ct_a[31] , \ct_a[30] , 
        \ct_a[29] , \ct_a[28] , \ct_a[27] , \ct_a[26] , \ct_a[25] , \ct_a[24] , 
        \ct_a[23] , \ct_a[22] , \ct_a[21] , \ct_a[20] , \ct_a[19] , \ct_a[18] , 
        \ct_a[17] , \ct_a[16] , \ct_a[15] , \ct_a[14] , \ct_a[13] , \ct_a[12] , 
        \ct_a[11] , \ct_a[10] , \ct_a[9] , \ct_a[8] , \ct_a[7] , \ct_a[6] , 
        \ct_a[5] , \ct_a[4] , \ct_a[3] , \ct_a[2] , \ct_a[1] , \ct_a[0] }), 
        .chainresponse(chainresponse), .crnw({\ct_rnw[1] , \ct_rnw[0] }), 
        .csize({\ct_size[3] , \ct_size[2] , \ct_size[1] , \ct_size[0] }), 
        .ctag({\ct_itag[9] , \ct_itag[8] , \ct_itag[7] , \ct_itag[6] , 
        \ct_itag[5] , \ct_itag[4] , \ct_itag[3] , \ct_itag[2] , \ct_itag[1] , 
        \ct_itag[0] }), .lock({\ct_lock[1] , \ct_lock[0] }), 
        .nchaincommandack(nchaincommandack), .nrouteack(nroute_ack), .rack(
        rt_ack), .routetxreq(routetx_req), .seq({\ct_seq[1] , \ct_seq[0] }), 
        .tag_h({\tag_h[4] , \tag_h[3] , \tag_h[2] , \tag_h[1] , \tag_h[0] }), 
        .tag_l({\tag_l[4] , \tag_l[3] , \tag_l[2] , \tag_l[1] , \tag_l[0] }), 
        .wd({\ct_wd[63] , \ct_wd[62] , \ct_wd[61] , \ct_wd[60] , \ct_wd[59] , 
        \ct_wd[58] , \ct_wd[57] , \ct_wd[56] , \ct_wd[55] , \ct_wd[54] , 
        \ct_wd[53] , \ct_wd[52] , \ct_wd[51] , \ct_wd[50] , \ct_wd[49] , 
        \ct_wd[48] , \ct_wd[47] , \ct_wd[46] , \ct_wd[45] , \ct_wd[44] , 
        \ct_wd[43] , \ct_wd[42] , \ct_wd[41] , \ct_wd[40] , \ct_wd[39] , 
        \ct_wd[38] , \ct_wd[37] , \ct_wd[36] , \ct_wd[35] , \ct_wd[34] , 
        \ct_wd[33] , \ct_wd[32] , \ct_wd[31] , \ct_wd[30] , \ct_wd[29] , 
        \ct_wd[28] , \ct_wd[27] , \ct_wd[26] , \ct_wd[25] , \ct_wd[24] , 
        \ct_wd[23] , \ct_wd[22] , \ct_wd[21] , \ct_wd[20] , \ct_wd[19] , 
        \ct_wd[18] , \ct_wd[17] , \ct_wd[16] , \ct_wd[15] , \ct_wd[14] , 
        \ct_wd[13] , \ct_wd[12] , \ct_wd[11] , \ct_wd[10] , \ct_wd[9] , 
        \ct_wd[8] , \ct_wd[7] , \ct_wd[6] , \ct_wd[5] , \ct_wd[4] , \ct_wd[3] , 
        \ct_wd[2] , \ct_wd[1] , \ct_wd[0] }), .cack(ct_ack), .cdefer(ct_defer), 
        .chaincommand(chaincommand), .cndefer(ct_slow), .cok(ct_ok), .err({
        \rt_err[1] , \rt_err[0] }), .nReset(nReset), .nchainresponseack(
        nchainresponseack), .rd({\rt_rd[63] , \rt_rd[62] , \rt_rd[61] , 
        \rt_rd[60] , \rt_rd[59] , \rt_rd[58] , \rt_rd[57] , \rt_rd[56] , 
        \rt_rd[55] , \rt_rd[54] , \rt_rd[53] , \rt_rd[52] , \rt_rd[51] , 
        \rt_rd[50] , \rt_rd[49] , \rt_rd[48] , \rt_rd[47] , \rt_rd[46] , 
        \rt_rd[45] , \rt_rd[44] , \rt_rd[43] , \rt_rd[42] , \rt_rd[41] , 
        \rt_rd[40] , \rt_rd[39] , \rt_rd[38] , \rt_rd[37] , \rt_rd[36] , 
        \rt_rd[35] , \rt_rd[34] , \rt_rd[33] , \rt_rd[32] , \rt_rd[31] , 
        \rt_rd[30] , \rt_rd[29] , \rt_rd[28] , \rt_rd[27] , \rt_rd[26] , 
        \rt_rd[25] , \rt_rd[24] , \rt_rd[23] , \rt_rd[22] , \rt_rd[21] , 
        \rt_rd[20] , \rt_rd[19] , \rt_rd[18] , \rt_rd[17] , \rt_rd[16] , 
        \rt_rd[15] , \rt_rd[14] , \rt_rd[13] , \rt_rd[12] , \rt_rd[11] , 
        \rt_rd[10] , \rt_rd[9] , \rt_rd[8] , \rt_rd[7] , \rt_rd[6] , 
        \rt_rd[5] , \rt_rd[4] , \rt_rd[3] , \rt_rd[2] , \rt_rd[1] , \rt_rd[0] 
        }), .route({\route[4] , 1'b0, 1'b0, \route[1] , \route[0] }), 
        .routetxack(routetx_ack) );
    t_adec_imem dec ( .e_h({SYNOPSYS_UNCONNECTED_1, \eh[1] , \eh[0] }), .e_l({
        \el[2] , \el[1] , \el[0] }), .r_h({\rh[2] , \rh[1] , 
        SYNOPSYS_UNCONNECTED_2}), .r_l({\rl[2] , \rl[1] , \rl[0] }), .e_dp(
        e_dp), .e_ip(e_ip), .e_tic(e_tic), .r_dp(r_dp), .r_ip(r_ip), .r_tic(
        r_tic), .tag_h({\tag_h[4] , \tag_h[3] , \tag_h[2] , \tag_h[1] , 
        \tag_h[0] }), .tag_l({\tag_l[4] , \tag_l[3] , \tag_l[2] , \tag_l[1] , 
        \tag_l[0] }) );
    resp_route_tx_imem rt ( .o({\route[4] , SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, \route[1] , \route[0] }), .rtxack(routetx_ack), 
        .e_h({1'b0, \eh[1] , \eh[0] }), .e_l({\el[2] , \el[1] , \el[0] }), 
        .noa(nroute_ack), .r_h({\rh[2] , \rh[1] , 1'b0}), .r_l({\rl[2] , 
        \rl[1] , \rl[0] }), .rtxreq(routetx_req) );
    inv_2 U1 ( .x(reset), .a(nReset) );
    cp2slave_imem chainif2slave ( .tc_seq({\ct_seq[1] , \ct_seq[0] }), 
        .tc_size({\ct_size[3] , \ct_size[2] , \ct_size[1] , \ct_size[0] }), 
        .tc_itag({\ct_itag[9] , \ct_itag[8] , \ct_itag[7] , \ct_itag[6] , 
        \ct_itag[5] , \ct_itag[4] , \ct_itag[3] , \ct_itag[2] , \ct_itag[1] , 
        \ct_itag[0] }), .tc_wd({\ct_wd[63] , \ct_wd[62] , \ct_wd[61] , 
        \ct_wd[60] , \ct_wd[59] , \ct_wd[58] , \ct_wd[57] , \ct_wd[56] , 
        \ct_wd[55] , \ct_wd[54] , \ct_wd[53] , \ct_wd[52] , \ct_wd[51] , 
        \ct_wd[50] , \ct_wd[49] , \ct_wd[48] , \ct_wd[47] , \ct_wd[46] , 
        \ct_wd[45] , \ct_wd[44] , \ct_wd[43] , \ct_wd[42] , \ct_wd[41] , 
        \ct_wd[40] , \ct_wd[39] , \ct_wd[38] , \ct_wd[37] , \ct_wd[36] , 
        \ct_wd[35] , \ct_wd[34] , \ct_wd[33] , \ct_wd[32] , \ct_wd[31] , 
        \ct_wd[30] , \ct_wd[29] , \ct_wd[28] , \ct_wd[27] , \ct_wd[26] , 
        \ct_wd[25] , \ct_wd[24] , \ct_wd[23] , \ct_wd[22] , \ct_wd[21] , 
        \ct_wd[20] , \ct_wd[19] , \ct_wd[18] , \ct_wd[17] , \ct_wd[16] , 
        \ct_wd[15] , \ct_wd[14] , \ct_wd[13] , \ct_wd[12] , \ct_wd[11] , 
        \ct_wd[10] , \ct_wd[9] , \ct_wd[8] , \ct_wd[7] , \ct_wd[6] , 
        \ct_wd[5] , \ct_wd[4] , \ct_wd[3] , \ct_wd[2] , \ct_wd[1] , \ct_wd[0] 
        }), .tc_lock({\ct_lock[1] , \ct_lock[0] }), .tc_a({\ct_a[63] , 
        \ct_a[62] , \ct_a[61] , \ct_a[60] , \ct_a[59] , \ct_a[58] , \ct_a[57] , 
        \ct_a[56] , \ct_a[55] , \ct_a[54] , \ct_a[53] , \ct_a[52] , \ct_a[51] , 
        \ct_a[50] , \ct_a[49] , \ct_a[48] , \ct_a[47] , \ct_a[46] , \ct_a[45] , 
        \ct_a[44] , \ct_a[43] , \ct_a[42] , \ct_a[41] , \ct_a[40] , \ct_a[39] , 
        \ct_a[38] , \ct_a[37] , \ct_a[36] , \ct_a[35] , \ct_a[34] , \ct_a[33] , 
        \ct_a[32] , \ct_a[31] , \ct_a[30] , \ct_a[29] , \ct_a[28] , \ct_a[27] , 
        \ct_a[26] , \ct_a[25] , \ct_a[24] , \ct_a[23] , \ct_a[22] , \ct_a[21] , 
        \ct_a[20] , \ct_a[19] , \ct_a[18] , \ct_a[17] , \ct_a[16] , \ct_a[15] , 
        \ct_a[14] , \ct_a[13] , \ct_a[12] , \ct_a[11] , \ct_a[10] , \ct_a[9] , 
        \ct_a[8] , \ct_a[7] , \ct_a[6] , \ct_a[5] , \ct_a[4] , \ct_a[3] , 
        \ct_a[2] , \ct_a[1] , \ct_a[0] }), .tc_rnw({\ct_rnw[1] , \ct_rnw[0] }), 
        .tc_ok(ct_ok), .tc_defer(ct_defer), .tc_slow(ct_slow), .tc_ack(ct_ack), 
        .req_in(sc_req), .st_i(sc_st), .we_i(sc_we), .mult_i(sc_mult), .adr_i(
        sc_adr), .dat_i(sc_dat), .seq_i(sc_seq), .sel_i({sc_sel[3], sc_sel[2], 
        sc_sel[1], SYNOPSYS_UNCONNECTED_5}), .ack_in(sc_ack), .tr_rd({
        \rt_rd[63] , \rt_rd[62] , \rt_rd[61] , \rt_rd[60] , \rt_rd[59] , 
        \rt_rd[58] , \rt_rd[57] , \rt_rd[56] , \rt_rd[55] , \rt_rd[54] , 
        \rt_rd[53] , \rt_rd[52] , \rt_rd[51] , \rt_rd[50] , \rt_rd[49] , 
        \rt_rd[48] , \rt_rd[47] , \rt_rd[46] , \rt_rd[45] , \rt_rd[44] , 
        \rt_rd[43] , \rt_rd[42] , \rt_rd[41] , \rt_rd[40] , \rt_rd[39] , 
        \rt_rd[38] , \rt_rd[37] , \rt_rd[36] , \rt_rd[35] , \rt_rd[34] , 
        \rt_rd[33] , \rt_rd[32] , \rt_rd[31] , \rt_rd[30] , \rt_rd[29] , 
        \rt_rd[28] , \rt_rd[27] , \rt_rd[26] , \rt_rd[25] , \rt_rd[24] , 
        \rt_rd[23] , \rt_rd[22] , \rt_rd[21] , \rt_rd[20] , \rt_rd[19] , 
        \rt_rd[18] , \rt_rd[17] , \rt_rd[16] , \rt_rd[15] , \rt_rd[14] , 
        \rt_rd[13] , \rt_rd[12] , \rt_rd[11] , \rt_rd[10] , \rt_rd[9] , 
        \rt_rd[8] , \rt_rd[7] , \rt_rd[6] , \rt_rd[5] , \rt_rd[4] , \rt_rd[3] , 
        \rt_rd[2] , \rt_rd[1] , \rt_rd[0] }), .tr_err({\rt_err[1] , 
        \rt_err[0] }), .tr_ack(rt_ack), .req_out(sr_req), .dat_o(sr_dat), 
        .err_o(sr_err), .rty_o(sr_rty), .acc_o(sr_acc), .sel_o(sr_sel), 
        .mult_o(sr_mult), .rt_o(sr_rt), .ack_out(sr_ack), .reset(reset) );
endmodule


module t_adec_dmem ( e_h, e_l, r_h, r_l, e_dp, e_ip, e_tic, r_dp, r_ip, r_tic, 
    tag_h, tag_l );
output [2:0] e_h;
output [2:0] e_l;
output [2:0] r_h;
output [2:0] r_l;
input  [2:0] e_dp;
input  [2:0] e_ip;
input  [2:0] e_tic;
input  [2:0] r_dp;
input  [2:0] r_ip;
input  [2:0] r_tic;
input  [4:0] tag_h;
input  [4:0] tag_l;
    wire \e_l[2] , \e_l[1] , \tag_h[4] , \e_l[0] ;
    assign e_h[2] = 1'b0;
    assign e_h[1] = \e_l[0] ;
    assign e_h[0] = \e_l[1] ;
    assign e_l[2] = \e_l[2] ;
    assign e_l[1] = \e_l[1] ;
    assign e_l[0] = \e_l[0] ;
    assign r_h[2] = \e_l[1] ;
    assign r_h[1] = \tag_h[4] ;
    assign r_h[0] = 1'b0;
    assign r_l[2] = \e_l[0] ;
    assign r_l[0] = \e_l[2] ;
    assign \tag_h[4]  = tag_h[4];
    or2_1 U3 ( .x(r_l[1]), .a(\e_l[0] ), .b(tag_h[3]) );
    buf_3 U6 ( .x(\e_l[0] ), .a(tag_h[2]) );
    or2_2 U7 ( .x(\e_l[1] ), .a(tag_h[3]), .b(\tag_h[4] ) );
    or2_2 U8 ( .x(\e_l[2] ), .a(\tag_h[4] ), .b(r_l[1]) );
endmodule


module chain_sendmux8_12 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/naa , \U1693/bdone , \U1693/net3 , 
        \U1693/drivemonitor , \U1693/net2 , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendmux8_13 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/naa , \U1693/bdone , \U1693/net3 , 
        \U1693/drivemonitor , \U1693/net2 , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendmux8_14 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/naa , \U1693/bdone , \U1693/net3 , 
        \U1693/drivemonitor , \U1693/net2 , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendmux8_15 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/naa , \U1693/bdone , \U1693/net3 , 
        \U1693/drivemonitor , \U1693/net2 , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendword_2 ( ctrlack, oh, ol, chainackff, ctrlreq, ih, il );
output [7:0] oh;
output [7:0] ol;
input  [31:0] ih;
input  [31:0] il;
input  chainackff, ctrlreq;
output ctrlack;
    wire \third_oh[7] , \third_oh[6] , \third_oh[5] , \third_oh[4] , 
        \third_oh[3] , \third_oh[2] , \third_oh[1] , \third_oh[0] , 
        \fourth_ol[7] , \fourth_ol[6] , \fourth_ol[5] , \fourth_ol[4] , 
        \fourth_ol[3] , \fourth_ol[2] , \fourth_ol[1] , \fourth_ol[0] , 
        \third_ol[7] , \third_ol[6] , \third_ol[5] , \third_ol[4] , 
        \third_ol[3] , \third_ol[2] , \third_ol[1] , \third_ol[0] , 
        \fourth_oh[7] , \fourth_oh[6] , \fourth_oh[5] , \fourth_oh[4] , 
        \fourth_oh[3] , \fourth_oh[2] , \fourth_oh[1] , \fourth_oh[0] , 
        \second_oh[7] , \second_oh[6] , \second_oh[5] , \second_oh[4] , 
        \second_oh[3] , \second_oh[2] , \second_oh[1] , \second_oh[0] , 
        \second_ol[7] , \second_ol[6] , \second_ol[5] , \second_ol[4] , 
        \second_ol[3] , \second_ol[2] , \second_ol[1] , \second_ol[0] , 
        \first_oh[7] , \first_oh[6] , \first_oh[5] , \first_oh[4] , 
        \first_oh[3] , \first_oh[2] , \first_oh[1] , \first_oh[0] , 
        \first_ol[7] , \first_ol[6] , \first_ol[5] , \first_ol[4] , 
        \first_ol[3] , \first_ol[2] , \first_ol[1] , \first_ol[0] , net44, 
        net51, net58, bctrlreq, \U309_0_/n5 , \U309_0_/n1 , \U309_0_/n2 , 
        \U309_0_/n3 , \U309_0_/n4 , \U309_1_/n5 , \U309_1_/n1 , \U309_1_/n2 , 
        \U309_1_/n3 , \U309_1_/n4 , \U309_2_/n5 , \U309_2_/n1 , \U309_2_/n2 , 
        \U309_2_/n3 , \U309_2_/n4 , \U309_3_/n5 , \U309_3_/n1 , \U309_3_/n2 , 
        \U309_3_/n3 , \U309_3_/n4 , \U309_4_/n5 , \U309_4_/n1 , \U309_4_/n2 , 
        \U309_4_/n3 , \U309_4_/n4 , \U309_5_/n5 , \U309_5_/n1 , \U309_5_/n2 , 
        \U309_5_/n3 , \U309_5_/n4 , \U309_6_/n5 , \U309_6_/n1 , \U309_6_/n2 , 
        \U309_6_/n3 , \U309_6_/n4 , \U309_7_/n5 , \U309_7_/n1 , \U309_7_/n2 , 
        \U309_7_/n3 , \U309_7_/n4 , \U310_0_/n5 , \U310_0_/n1 , \U310_0_/n2 , 
        \U310_0_/n3 , \U310_0_/n4 , \U310_1_/n5 , \U310_1_/n1 , \U310_1_/n2 , 
        \U310_1_/n3 , \U310_1_/n4 , \U310_2_/n5 , \U310_2_/n1 , \U310_2_/n2 , 
        \U310_2_/n3 , \U310_2_/n4 , \U310_3_/n5 , \U310_3_/n1 , \U310_3_/n2 , 
        \U310_3_/n3 , \U310_3_/n4 , \U310_4_/n5 , \U310_4_/n1 , \U310_4_/n2 , 
        \U310_4_/n3 , \U310_4_/n4 , \U310_5_/n5 , \U310_5_/n1 , \U310_5_/n2 , 
        \U310_5_/n3 , \U310_5_/n4 , \U310_6_/n5 , \U310_6_/n1 , \U310_6_/n2 , 
        \U310_6_/n3 , \U310_6_/n4 , \U310_7_/n5 , \U310_7_/n1 , \U310_7_/n2 , 
        \U310_7_/n3 , \U310_7_/n4 ;
    chain_sendmux8_14 I4 ( .ctrlack(ctrlack), .oh({\fourth_oh[7] , 
        \fourth_oh[6] , \fourth_oh[5] , \fourth_oh[4] , \fourth_oh[3] , 
        \fourth_oh[2] , \fourth_oh[1] , \fourth_oh[0] }), .ol({\fourth_ol[7] , 
        \fourth_ol[6] , \fourth_ol[5] , \fourth_ol[4] , \fourth_ol[3] , 
        \fourth_ol[2] , \fourth_ol[1] , \fourth_ol[0] }), .i_h(ih[7:0]), .i_l(
        il[7:0]), .ctrlreq(net44), .oa(chainackff) );
    chain_sendmux8_13 I3 ( .ctrlack(net44), .oh({\third_oh[7] , \third_oh[6] , 
        \third_oh[5] , \third_oh[4] , \third_oh[3] , \third_oh[2] , 
        \third_oh[1] , \third_oh[0] }), .ol({\third_ol[7] , \third_ol[6] , 
        \third_ol[5] , \third_ol[4] , \third_ol[3] , \third_ol[2] , 
        \third_ol[1] , \third_ol[0] }), .i_h(ih[15:8]), .i_l(il[15:8]), 
        .ctrlreq(net51), .oa(chainackff) );
    chain_sendmux8_12 I2 ( .ctrlack(net51), .oh({\second_oh[7] , 
        \second_oh[6] , \second_oh[5] , \second_oh[4] , \second_oh[3] , 
        \second_oh[2] , \second_oh[1] , \second_oh[0] }), .ol({\second_ol[7] , 
        \second_ol[6] , \second_ol[5] , \second_ol[4] , \second_ol[3] , 
        \second_ol[2] , \second_ol[1] , \second_ol[0] }), .i_h(ih[23:16]), 
        .i_l(il[23:16]), .ctrlreq(net58), .oa(chainackff) );
    chain_sendmux8_15 U320 ( .ctrlack(net58), .oh({\first_oh[7] , 
        \first_oh[6] , \first_oh[5] , \first_oh[4] , \first_oh[3] , 
        \first_oh[2] , \first_oh[1] , \first_oh[0] }), .ol({\first_ol[7] , 
        \first_ol[6] , \first_ol[5] , \first_ol[4] , \first_ol[3] , 
        \first_ol[2] , \first_ol[1] , \first_ol[0] }), .i_h(ih[31:24]), .i_l(
        il[31:24]), .ctrlreq(bctrlreq), .oa(chainackff) );
    buf_2 \U328/U7  ( .x(bctrlreq), .a(ctrlreq) );
    and4_2 \U309_0_/U24  ( .x(\U309_0_/n5 ), .a(\U309_0_/n1 ), .b(\U309_0_/n2 
        ), .c(\U309_0_/n3 ), .d(\U309_0_/n4 ) );
    inv_1 \U309_0_/U1  ( .x(\U309_0_/n1 ), .a(\fourth_oh[0] ) );
    inv_1 \U309_0_/U2  ( .x(\U309_0_/n2 ), .a(\third_oh[0] ) );
    inv_1 \U309_0_/U3  ( .x(\U309_0_/n3 ), .a(\second_oh[0] ) );
    inv_1 \U309_0_/U4  ( .x(\U309_0_/n4 ), .a(\first_oh[0] ) );
    inv_4 \U309_0_/U5  ( .x(oh[0]), .a(\U309_0_/n5 ) );
    and4_2 \U309_1_/U24  ( .x(\U309_1_/n5 ), .a(\U309_1_/n1 ), .b(\U309_1_/n2 
        ), .c(\U309_1_/n3 ), .d(\U309_1_/n4 ) );
    inv_1 \U309_1_/U1  ( .x(\U309_1_/n1 ), .a(\fourth_oh[1] ) );
    inv_1 \U309_1_/U2  ( .x(\U309_1_/n2 ), .a(\third_oh[1] ) );
    inv_1 \U309_1_/U3  ( .x(\U309_1_/n3 ), .a(\second_oh[1] ) );
    inv_1 \U309_1_/U4  ( .x(\U309_1_/n4 ), .a(\first_oh[1] ) );
    inv_4 \U309_1_/U5  ( .x(oh[1]), .a(\U309_1_/n5 ) );
    and4_2 \U309_2_/U24  ( .x(\U309_2_/n5 ), .a(\U309_2_/n1 ), .b(\U309_2_/n2 
        ), .c(\U309_2_/n3 ), .d(\U309_2_/n4 ) );
    inv_1 \U309_2_/U1  ( .x(\U309_2_/n1 ), .a(\fourth_oh[2] ) );
    inv_1 \U309_2_/U2  ( .x(\U309_2_/n2 ), .a(\third_oh[2] ) );
    inv_1 \U309_2_/U3  ( .x(\U309_2_/n3 ), .a(\second_oh[2] ) );
    inv_1 \U309_2_/U4  ( .x(\U309_2_/n4 ), .a(\first_oh[2] ) );
    inv_4 \U309_2_/U5  ( .x(oh[2]), .a(\U309_2_/n5 ) );
    and4_2 \U309_3_/U24  ( .x(\U309_3_/n5 ), .a(\U309_3_/n1 ), .b(\U309_3_/n2 
        ), .c(\U309_3_/n3 ), .d(\U309_3_/n4 ) );
    inv_1 \U309_3_/U1  ( .x(\U309_3_/n1 ), .a(\fourth_oh[3] ) );
    inv_1 \U309_3_/U2  ( .x(\U309_3_/n2 ), .a(\third_oh[3] ) );
    inv_1 \U309_3_/U3  ( .x(\U309_3_/n3 ), .a(\second_oh[3] ) );
    inv_1 \U309_3_/U4  ( .x(\U309_3_/n4 ), .a(\first_oh[3] ) );
    inv_4 \U309_3_/U5  ( .x(oh[3]), .a(\U309_3_/n5 ) );
    and4_2 \U309_4_/U24  ( .x(\U309_4_/n5 ), .a(\U309_4_/n1 ), .b(\U309_4_/n2 
        ), .c(\U309_4_/n3 ), .d(\U309_4_/n4 ) );
    inv_1 \U309_4_/U1  ( .x(\U309_4_/n1 ), .a(\fourth_oh[4] ) );
    inv_1 \U309_4_/U2  ( .x(\U309_4_/n2 ), .a(\third_oh[4] ) );
    inv_1 \U309_4_/U3  ( .x(\U309_4_/n3 ), .a(\second_oh[4] ) );
    inv_1 \U309_4_/U4  ( .x(\U309_4_/n4 ), .a(\first_oh[4] ) );
    inv_4 \U309_4_/U5  ( .x(oh[4]), .a(\U309_4_/n5 ) );
    and4_2 \U309_5_/U24  ( .x(\U309_5_/n5 ), .a(\U309_5_/n1 ), .b(\U309_5_/n2 
        ), .c(\U309_5_/n3 ), .d(\U309_5_/n4 ) );
    inv_1 \U309_5_/U1  ( .x(\U309_5_/n1 ), .a(\fourth_oh[5] ) );
    inv_1 \U309_5_/U2  ( .x(\U309_5_/n2 ), .a(\third_oh[5] ) );
    inv_1 \U309_5_/U3  ( .x(\U309_5_/n3 ), .a(\second_oh[5] ) );
    inv_1 \U309_5_/U4  ( .x(\U309_5_/n4 ), .a(\first_oh[5] ) );
    inv_4 \U309_5_/U5  ( .x(oh[5]), .a(\U309_5_/n5 ) );
    and4_2 \U309_6_/U24  ( .x(\U309_6_/n5 ), .a(\U309_6_/n1 ), .b(\U309_6_/n2 
        ), .c(\U309_6_/n3 ), .d(\U309_6_/n4 ) );
    inv_1 \U309_6_/U1  ( .x(\U309_6_/n1 ), .a(\fourth_oh[6] ) );
    inv_1 \U309_6_/U2  ( .x(\U309_6_/n2 ), .a(\third_oh[6] ) );
    inv_1 \U309_6_/U3  ( .x(\U309_6_/n3 ), .a(\second_oh[6] ) );
    inv_1 \U309_6_/U4  ( .x(\U309_6_/n4 ), .a(\first_oh[6] ) );
    inv_4 \U309_6_/U5  ( .x(oh[6]), .a(\U309_6_/n5 ) );
    and4_2 \U309_7_/U24  ( .x(\U309_7_/n5 ), .a(\U309_7_/n1 ), .b(\U309_7_/n2 
        ), .c(\U309_7_/n3 ), .d(\U309_7_/n4 ) );
    inv_1 \U309_7_/U1  ( .x(\U309_7_/n1 ), .a(\fourth_oh[7] ) );
    inv_1 \U309_7_/U2  ( .x(\U309_7_/n2 ), .a(\third_oh[7] ) );
    inv_1 \U309_7_/U3  ( .x(\U309_7_/n3 ), .a(\second_oh[7] ) );
    inv_1 \U309_7_/U4  ( .x(\U309_7_/n4 ), .a(\first_oh[7] ) );
    inv_4 \U309_7_/U5  ( .x(oh[7]), .a(\U309_7_/n5 ) );
    and4_2 \U310_0_/U24  ( .x(\U310_0_/n5 ), .a(\U310_0_/n1 ), .b(\U310_0_/n2 
        ), .c(\U310_0_/n3 ), .d(\U310_0_/n4 ) );
    inv_1 \U310_0_/U1  ( .x(\U310_0_/n1 ), .a(\fourth_ol[0] ) );
    inv_1 \U310_0_/U2  ( .x(\U310_0_/n2 ), .a(\third_ol[0] ) );
    inv_1 \U310_0_/U3  ( .x(\U310_0_/n3 ), .a(\second_ol[0] ) );
    inv_1 \U310_0_/U4  ( .x(\U310_0_/n4 ), .a(\first_ol[0] ) );
    inv_4 \U310_0_/U5  ( .x(ol[0]), .a(\U310_0_/n5 ) );
    and4_2 \U310_1_/U24  ( .x(\U310_1_/n5 ), .a(\U310_1_/n1 ), .b(\U310_1_/n2 
        ), .c(\U310_1_/n3 ), .d(\U310_1_/n4 ) );
    inv_1 \U310_1_/U1  ( .x(\U310_1_/n1 ), .a(\fourth_ol[1] ) );
    inv_1 \U310_1_/U2  ( .x(\U310_1_/n2 ), .a(\third_ol[1] ) );
    inv_1 \U310_1_/U3  ( .x(\U310_1_/n3 ), .a(\second_ol[1] ) );
    inv_1 \U310_1_/U4  ( .x(\U310_1_/n4 ), .a(\first_ol[1] ) );
    inv_4 \U310_1_/U5  ( .x(ol[1]), .a(\U310_1_/n5 ) );
    and4_2 \U310_2_/U24  ( .x(\U310_2_/n5 ), .a(\U310_2_/n1 ), .b(\U310_2_/n2 
        ), .c(\U310_2_/n3 ), .d(\U310_2_/n4 ) );
    inv_1 \U310_2_/U1  ( .x(\U310_2_/n1 ), .a(\fourth_ol[2] ) );
    inv_1 \U310_2_/U2  ( .x(\U310_2_/n2 ), .a(\third_ol[2] ) );
    inv_1 \U310_2_/U3  ( .x(\U310_2_/n3 ), .a(\second_ol[2] ) );
    inv_1 \U310_2_/U4  ( .x(\U310_2_/n4 ), .a(\first_ol[2] ) );
    inv_4 \U310_2_/U5  ( .x(ol[2]), .a(\U310_2_/n5 ) );
    and4_2 \U310_3_/U24  ( .x(\U310_3_/n5 ), .a(\U310_3_/n1 ), .b(\U310_3_/n2 
        ), .c(\U310_3_/n3 ), .d(\U310_3_/n4 ) );
    inv_1 \U310_3_/U1  ( .x(\U310_3_/n1 ), .a(\fourth_ol[3] ) );
    inv_1 \U310_3_/U2  ( .x(\U310_3_/n2 ), .a(\third_ol[3] ) );
    inv_1 \U310_3_/U3  ( .x(\U310_3_/n3 ), .a(\second_ol[3] ) );
    inv_1 \U310_3_/U4  ( .x(\U310_3_/n4 ), .a(\first_ol[3] ) );
    inv_4 \U310_3_/U5  ( .x(ol[3]), .a(\U310_3_/n5 ) );
    and4_2 \U310_4_/U24  ( .x(\U310_4_/n5 ), .a(\U310_4_/n1 ), .b(\U310_4_/n2 
        ), .c(\U310_4_/n3 ), .d(\U310_4_/n4 ) );
    inv_1 \U310_4_/U1  ( .x(\U310_4_/n1 ), .a(\fourth_ol[4] ) );
    inv_1 \U310_4_/U2  ( .x(\U310_4_/n2 ), .a(\third_ol[4] ) );
    inv_1 \U310_4_/U3  ( .x(\U310_4_/n3 ), .a(\second_ol[4] ) );
    inv_1 \U310_4_/U4  ( .x(\U310_4_/n4 ), .a(\first_ol[4] ) );
    inv_4 \U310_4_/U5  ( .x(ol[4]), .a(\U310_4_/n5 ) );
    and4_2 \U310_5_/U24  ( .x(\U310_5_/n5 ), .a(\U310_5_/n1 ), .b(\U310_5_/n2 
        ), .c(\U310_5_/n3 ), .d(\U310_5_/n4 ) );
    inv_1 \U310_5_/U1  ( .x(\U310_5_/n1 ), .a(\fourth_ol[5] ) );
    inv_1 \U310_5_/U2  ( .x(\U310_5_/n2 ), .a(\third_ol[5] ) );
    inv_1 \U310_5_/U3  ( .x(\U310_5_/n3 ), .a(\second_ol[5] ) );
    inv_1 \U310_5_/U4  ( .x(\U310_5_/n4 ), .a(\first_ol[5] ) );
    inv_4 \U310_5_/U5  ( .x(ol[5]), .a(\U310_5_/n5 ) );
    and4_2 \U310_6_/U24  ( .x(\U310_6_/n5 ), .a(\U310_6_/n1 ), .b(\U310_6_/n2 
        ), .c(\U310_6_/n3 ), .d(\U310_6_/n4 ) );
    inv_1 \U310_6_/U1  ( .x(\U310_6_/n1 ), .a(\fourth_ol[6] ) );
    inv_1 \U310_6_/U2  ( .x(\U310_6_/n2 ), .a(\third_ol[6] ) );
    inv_1 \U310_6_/U3  ( .x(\U310_6_/n3 ), .a(\second_ol[6] ) );
    inv_1 \U310_6_/U4  ( .x(\U310_6_/n4 ), .a(\first_ol[6] ) );
    inv_4 \U310_6_/U5  ( .x(ol[6]), .a(\U310_6_/n5 ) );
    and4_2 \U310_7_/U24  ( .x(\U310_7_/n5 ), .a(\U310_7_/n1 ), .b(\U310_7_/n2 
        ), .c(\U310_7_/n3 ), .d(\U310_7_/n4 ) );
    inv_1 \U310_7_/U1  ( .x(\U310_7_/n1 ), .a(\fourth_ol[7] ) );
    inv_1 \U310_7_/U2  ( .x(\U310_7_/n2 ), .a(\third_ol[7] ) );
    inv_1 \U310_7_/U3  ( .x(\U310_7_/n3 ), .a(\second_ol[7] ) );
    inv_1 \U310_7_/U4  ( .x(\U310_7_/n4 ), .a(\first_ol[7] ) );
    inv_4 \U310_7_/U5  ( .x(ol[7]), .a(\U310_7_/n5 ) );
endmodule


module chain_selement_ga_65 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_trhdr_2 ( chainff_ack, chainh, chainl, eop, hdrack, normal_ack, 
    notify_ack, read_req, routereq, chain_ff_h, chainack, chainff_l, eopack, 
    err, nReset, normal_response, notify_accept, notify_defer, rcol_h, rcol_l, 
    read_ack, rnw_h, rnw_l, routeack, rsize_h, rsize_l, rtag_h, rtag_l );
output [7:0] chainh;
output [7:0] chainl;
input  [7:0] chain_ff_h;
input  [7:0] chainff_l;
input  [1:0] err;
input  [2:0] rcol_h;
input  [2:0] rcol_l;
input  [1:0] rsize_h;
input  [1:0] rsize_l;
input  [4:0] rtag_h;
input  [4:0] rtag_l;
input  chainack, eopack, nReset, normal_response, notify_accept, notify_defer, 
    read_ack, rnw_h, rnw_l, routeack;
output chainff_ack, eop, hdrack, normal_ack, notify_ack, read_req, routereq;
    wire \net334[0] , \net334[1] , \net334[2] , \net334[4] , \net334[6] , 
        \net334[7] , \net413[0] , \net413[1] , \net413[2] , \net413[3] , 
        \net413[4] , \net413[5] , \net413[6] , \net413[7] , \net413[8] , 
        \net413[9] , \net413[10] , \net413[11] , \net413[12] , \net413[13] , 
        \net413[14] , \net413[15] , \net284[0] , \net284[1] , \net284[2] , 
        \net284[3] , \net284[4] , \net284[5] , \net284[6] , \net284[7] , 
        \net288[0] , \net288[1] , \net288[2] , \net288[3] , \net288[4] , 
        \net288[5] , \net288[6] , \net288[7] , \net343[0] , \net343[1] , 
        \net343[2] , \net343[3] , \net343[5] , \net343[6] , \net343[7] , 
        \hdr[17] , \hdr[16] , \hdr[1] , \hdr[0] , \drive_h[1] , \drive_h[0] , 
        \drive_l[1] , \drive_l[0] , done_write, dowrite, done_eop, ctrl_cd, 
        done_read, done_hdr, done_defer, net321, net362, net359, done_accept, 
        net332, net337, net340, done_pl, net364, donotify, net383, net0230, 
        net407, \U319/U21/U1/loop , \U323/U21/U1/loop , \U320/U21/U1/loop , 
        \U321/U21/U1/loop , \U322/U21/U1/loop , \U311/U28/Z , \U311/U32/Z , 
        \U311/U20/Z , \U311/U29/Z , \U311/U25/Z , \U311/U33/Z , \U311/U21/Z , 
        \U311/U26/Z , \U311/U34/Z , \U311/U30/Z , \U311/U19/Z , \U311/U27/Z , 
        \U311/U35/Z , \U311/U31/Z , \U311/nz[0] , \U311/nz[1] , \U311/x[1] , 
        \U311/y[3] , \U311/y[2] , \U311/x[7] , \U311/x[6] , \U311/x[4] , 
        \U311/y[1] , \U311/x[3] , \U311/x[2] , \U311/y[0] , \U311/x[5] , 
        \U311/x[0] , \U151/Z , \U210/naa , \U210/bdone , \U210/net3 , 
        \U210/drivemonitor , \U210/net2 , \U210/U1702/Z , \I0/naa , \I0/bdone , 
        \I0/net3 , \I0/drivemonitor , \I0/net2 , \I0/U1702/Z ;
    chain_selement_ga_65 U215 ( .Aa(done_eop), .Br(eop), .Ar(done_pl), .Ba(
        eopack) );
    nor2_1 \U308_0_/U5  ( .x(\net413[15] ), .a(\hdr[16] ), .b(\hdr[0] ) );
    nor2_1 \U308_1_/U5  ( .x(\net413[14] ), .a(\hdr[17] ), .b(\hdr[1] ) );
    nor2_1 \U308_2_/U5  ( .x(\net413[13] ), .a(1'b0), .b(routereq) );
    nor2_1 \U308_3_/U5  ( .x(\net413[12] ), .a(routereq), .b(1'b0) );
    nor2_1 \U308_4_/U5  ( .x(\net413[11] ), .a(1'b0), .b(routereq) );
    nor2_1 \U308_5_/U5  ( .x(\net413[10] ), .a(rnw_h), .b(rnw_l) );
    nor2_1 \U308_6_/U5  ( .x(\net413[9] ), .a(rsize_h[0]), .b(rsize_l[0]) );
    nor2_1 \U308_7_/U5  ( .x(\net413[8] ), .a(rsize_h[1]), .b(rsize_l[1]) );
    nor2_1 \U308_8_/U5  ( .x(\net413[7] ), .a(rtag_h[0]), .b(rtag_l[0]) );
    nor2_1 \U308_9_/U5  ( .x(\net413[6] ), .a(rtag_h[1]), .b(rtag_l[1]) );
    nor2_1 \U308_10_/U5  ( .x(\net413[5] ), .a(rtag_h[2]), .b(rtag_l[2]) );
    nor2_1 \U308_11_/U5  ( .x(\net413[4] ), .a(rtag_h[3]), .b(rtag_l[3]) );
    nor2_1 \U308_12_/U5  ( .x(\net413[3] ), .a(rtag_h[4]), .b(rtag_l[4]) );
    nor2_1 \U308_13_/U5  ( .x(\net413[2] ), .a(rcol_h[0]), .b(rcol_l[0]) );
    nor2_1 \U308_14_/U5  ( .x(\net413[1] ), .a(rcol_h[1]), .b(rcol_l[1]) );
    nor2_1 \U308_15_/U5  ( .x(\net413[0] ), .a(rcol_h[2]), .b(rcol_l[2]) );
    or3_1 \U257/U12  ( .x(net364), .a(donotify), .b(dowrite), .c(read_ack) );
    or3_1 \U297/U12  ( .x(net383), .a(done_defer), .b(done_write), .c(
        done_read) );
    and2_2 \U237/U8  ( .x(\hdr[1] ), .a(nReset), .b(normal_response) );
    and2_1 \U307_0_/U8  ( .x(\net343[7] ), .a(\drive_l[0] ), .b(\hdr[0] ) );
    and2_1 \U307_1_/U8  ( .x(\net343[6] ), .a(\drive_l[0] ), .b(\hdr[1] ) );
    and2_1 \U307_2_/U8  ( .x(\net343[5] ), .a(\drive_l[0] ), .b(routereq) );
    and2_1 \U307_4_/U8  ( .x(\net343[3] ), .a(\drive_l[0] ), .b(routereq) );
    and2_1 \U307_5_/U8  ( .x(\net343[2] ), .a(\drive_l[0] ), .b(rnw_l) );
    and2_1 \U307_6_/U8  ( .x(\net343[1] ), .a(\drive_l[0] ), .b(rsize_l[0]) );
    and2_1 \U307_7_/U8  ( .x(\net343[0] ), .a(\drive_l[0] ), .b(rsize_l[1]) );
    and2_1 \U235/U8  ( .x(net340), .a(err[1]), .b(nReset) );
    and2_1 \U236/U8  ( .x(net337), .a(nReset), .b(err[0]) );
    and2_1 \U306_0_/U8  ( .x(\net334[7] ), .a(\hdr[16] ), .b(\drive_l[1] ) );
    and2_1 \U306_1_/U8  ( .x(\net334[6] ), .a(\hdr[17] ), .b(\drive_l[1] ) );
    and2_1 \U306_3_/U8  ( .x(\net334[4] ), .a(routereq), .b(\drive_l[1] ) );
    and2_1 \U306_5_/U8  ( .x(\net334[2] ), .a(rnw_h), .b(\drive_l[1] ) );
    and2_1 \U306_6_/U8  ( .x(\net334[1] ), .a(rsize_h[0]), .b(\drive_l[1] ) );
    and2_1 \U306_7_/U8  ( .x(\net334[0] ), .a(rsize_h[1]), .b(\drive_l[1] ) );
    and2_1 \I1_0_/U8  ( .x(\net284[7] ), .a(rtag_h[0]), .b(\drive_h[1] ) );
    and2_1 \I1_1_/U8  ( .x(\net284[6] ), .a(rtag_h[1]), .b(\drive_h[1] ) );
    and2_1 \I1_2_/U8  ( .x(\net284[5] ), .a(rtag_h[2]), .b(\drive_h[1] ) );
    and2_1 \I1_3_/U8  ( .x(\net284[4] ), .a(rtag_h[3]), .b(\drive_h[1] ) );
    and2_1 \I1_4_/U8  ( .x(\net284[3] ), .a(rtag_h[4]), .b(\drive_h[1] ) );
    and2_1 \I1_5_/U8  ( .x(\net284[2] ), .a(rcol_h[0]), .b(\drive_h[1] ) );
    and2_1 \I1_6_/U8  ( .x(\net284[1] ), .a(rcol_h[1]), .b(\drive_h[1] ) );
    and2_1 \I1_7_/U8  ( .x(\net284[0] ), .a(rcol_h[2]), .b(\drive_h[1] ) );
    and2_1 \I2_0_/U8  ( .x(\net288[7] ), .a(\drive_h[0] ), .b(rtag_l[0]) );
    and2_1 \I2_1_/U8  ( .x(\net288[6] ), .a(\drive_h[0] ), .b(rtag_l[1]) );
    and2_1 \I2_2_/U8  ( .x(\net288[5] ), .a(\drive_h[0] ), .b(rtag_l[2]) );
    and2_1 \I2_3_/U8  ( .x(\net288[4] ), .a(\drive_h[0] ), .b(rtag_l[3]) );
    and2_1 \I2_4_/U8  ( .x(\net288[3] ), .a(\drive_h[0] ), .b(rtag_l[4]) );
    and2_1 \I2_5_/U8  ( .x(\net288[2] ), .a(\drive_h[0] ), .b(rcol_l[0]) );
    and2_1 \I2_6_/U8  ( .x(\net288[1] ), .a(\drive_h[0] ), .b(rcol_l[1]) );
    and2_1 \I2_7_/U8  ( .x(\net288[0] ), .a(\drive_h[0] ), .b(rcol_l[2]) );
    inv_1 \U318/U3  ( .x(net332), .a(routereq) );
    or2_4 \U255/U12  ( .x(notify_ack), .a(done_accept), .b(done_defer) );
    or2_4 \U228/U12  ( .x(\hdr[17] ), .a(notify_defer), .b(notify_accept) );
    or2_4 \U204/U12  ( .x(net321), .a(net359), .b(net362) );
    or2_4 \U221/U12  ( .x(\hdr[16] ), .a(net359), .b(notify_defer) );
    or2_4 \U252/U12  ( .x(normal_ack), .a(done_write), .b(done_read) );
    or2_4 \U280/U12  ( .x(\hdr[0] ), .a(net362), .b(notify_accept) );
    or2_4 \U317/U12  ( .x(routereq), .a(\hdr[17] ), .b(net321) );
    or3_4 \U309_0_/U12  ( .x(chainh[0]), .a(\net334[7] ), .b(\net284[7] ), .c(
        chain_ff_h[0]) );
    or3_4 \U309_1_/U12  ( .x(chainh[1]), .a(\net334[6] ), .b(\net284[6] ), .c(
        chain_ff_h[1]) );
    or3_4 \U309_3_/U12  ( .x(chainh[3]), .a(\net334[4] ), .b(\net284[4] ), .c(
        chain_ff_h[3]) );
    or3_4 \U309_5_/U12  ( .x(chainh[5]), .a(\net334[2] ), .b(\net284[2] ), .c(
        chain_ff_h[5]) );
    or3_4 \U309_6_/U12  ( .x(chainh[6]), .a(\net334[1] ), .b(\net284[1] ), .c(
        chain_ff_h[6]) );
    or3_4 \U309_7_/U12  ( .x(chainh[7]), .a(\net334[0] ), .b(\net284[0] ), .c(
        chain_ff_h[7]) );
    or3_4 \U310_0_/U12  ( .x(chainl[0]), .a(\net343[7] ), .b(\net288[7] ), .c(
        chainff_l[0]) );
    or3_4 \U310_1_/U12  ( .x(chainl[1]), .a(\net343[6] ), .b(\net288[6] ), .c(
        chainff_l[1]) );
    or3_4 \U310_2_/U12  ( .x(chainl[2]), .a(\net343[5] ), .b(\net288[5] ), .c(
        chainff_l[2]) );
    or3_4 \U310_4_/U12  ( .x(chainl[4]), .a(\net343[3] ), .b(\net288[3] ), .c(
        chainff_l[4]) );
    or3_4 \U310_5_/U12  ( .x(chainl[5]), .a(\net343[2] ), .b(\net288[2] ), .c(
        chainff_l[5]) );
    or3_4 \U310_6_/U12  ( .x(chainl[6]), .a(\net343[1] ), .b(\net288[1] ), .c(
        chainff_l[6]) );
    or3_4 \U310_7_/U12  ( .x(chainl[7]), .a(\net343[0] ), .b(\net288[0] ), .c(
        chainff_l[7]) );
    ao222_1 \U311/U37/U18/U1/U1  ( .x(ctrl_cd), .a(\U311/nz[0] ), .b(
        \U311/nz[1] ), .c(\U311/nz[0] ), .d(ctrl_cd), .e(\U311/nz[1] ), .f(
        ctrl_cd) );
    aoi222_1 \U311/U28/U30/U1  ( .x(\U311/x[3] ), .a(\net413[8] ), .b(
        \net413[9] ), .c(\net413[8] ), .d(\U311/U28/Z ), .e(\net413[9] ), .f(
        \U311/U28/Z ) );
    inv_1 \U311/U28/U30/Uinv  ( .x(\U311/U28/Z ), .a(\U311/x[3] ) );
    aoi222_1 \U311/U32/U30/U1  ( .x(\U311/x[0] ), .a(\net413[14] ), .b(
        \net413[15] ), .c(\net413[14] ), .d(\U311/U32/Z ), .e(\net413[15] ), 
        .f(\U311/U32/Z ) );
    inv_1 \U311/U32/U30/Uinv  ( .x(\U311/U32/Z ), .a(\U311/x[0] ) );
    aoi222_1 \U311/U20/U30/U1  ( .x(\U311/x[5] ), .a(\net413[4] ), .b(
        \net413[5] ), .c(\net413[4] ), .d(\U311/U20/Z ), .e(\net413[5] ), .f(
        \U311/U20/Z ) );
    inv_1 \U311/U20/U30/Uinv  ( .x(\U311/U20/Z ), .a(\U311/x[5] ) );
    aoi222_1 \U311/U29/U30/U1  ( .x(\U311/x[2] ), .a(\net413[10] ), .b(
        \net413[11] ), .c(\net413[10] ), .d(\U311/U29/Z ), .e(\net413[11] ), 
        .f(\U311/U29/Z ) );
    inv_1 \U311/U29/U30/Uinv  ( .x(\U311/U29/Z ), .a(\U311/x[2] ) );
    aoi222_1 \U311/U25/U30/U1  ( .x(\U311/x[7] ), .a(\net413[0] ), .b(
        \net413[1] ), .c(\net413[0] ), .d(\U311/U25/Z ), .e(\net413[1] ), .f(
        \U311/U25/Z ) );
    inv_1 \U311/U25/U30/Uinv  ( .x(\U311/U25/Z ), .a(\U311/x[7] ) );
    aoi222_1 \U311/U33/U30/U1  ( .x(\U311/y[0] ), .a(\U311/x[1] ), .b(
        \U311/x[0] ), .c(\U311/x[1] ), .d(\U311/U33/Z ), .e(\U311/x[0] ), .f(
        \U311/U33/Z ) );
    inv_1 \U311/U33/U30/Uinv  ( .x(\U311/U33/Z ), .a(\U311/y[0] ) );
    aoi222_1 \U311/U21/U30/U1  ( .x(\U311/y[2] ), .a(\U311/x[5] ), .b(
        \U311/x[4] ), .c(\U311/x[5] ), .d(\U311/U21/Z ), .e(\U311/x[4] ), .f(
        \U311/U21/Z ) );
    inv_1 \U311/U21/U30/Uinv  ( .x(\U311/U21/Z ), .a(\U311/y[2] ) );
    aoi222_1 \U311/U26/U30/U1  ( .x(\U311/x[6] ), .a(\net413[2] ), .b(
        \net413[3] ), .c(\net413[2] ), .d(\U311/U26/Z ), .e(\net413[3] ), .f(
        \U311/U26/Z ) );
    inv_1 \U311/U26/U30/Uinv  ( .x(\U311/U26/Z ), .a(\U311/x[6] ) );
    aoi222_1 \U311/U34/U30/U1  ( .x(\U311/nz[0] ), .a(\U311/y[1] ), .b(
        \U311/y[0] ), .c(\U311/y[1] ), .d(\U311/U34/Z ), .e(\U311/y[0] ), .f(
        \U311/U34/Z ) );
    inv_1 \U311/U34/U30/Uinv  ( .x(\U311/U34/Z ), .a(\U311/nz[0] ) );
    aoi222_1 \U311/U30/U30/U1  ( .x(\U311/y[1] ), .a(\U311/x[3] ), .b(
        \U311/x[2] ), .c(\U311/x[3] ), .d(\U311/U30/Z ), .e(\U311/x[2] ), .f(
        \U311/U30/Z ) );
    inv_1 \U311/U30/U30/Uinv  ( .x(\U311/U30/Z ), .a(\U311/y[1] ) );
    aoi222_1 \U311/U19/U30/U1  ( .x(\U311/x[4] ), .a(\net413[6] ), .b(
        \net413[7] ), .c(\net413[6] ), .d(\U311/U19/Z ), .e(\net413[7] ), .f(
        \U311/U19/Z ) );
    inv_1 \U311/U19/U30/Uinv  ( .x(\U311/U19/Z ), .a(\U311/x[4] ) );
    aoi222_1 \U311/U27/U30/U1  ( .x(\U311/y[3] ), .a(\U311/x[7] ), .b(
        \U311/x[6] ), .c(\U311/x[7] ), .d(\U311/U27/Z ), .e(\U311/x[6] ), .f(
        \U311/U27/Z ) );
    inv_1 \U311/U27/U30/Uinv  ( .x(\U311/U27/Z ), .a(\U311/y[3] ) );
    aoi222_1 \U311/U35/U30/U1  ( .x(\U311/nz[1] ), .a(\U311/y[3] ), .b(
        \U311/y[2] ), .c(\U311/y[3] ), .d(\U311/U35/Z ), .e(\U311/y[2] ), .f(
        \U311/U35/Z ) );
    inv_1 \U311/U35/U30/Uinv  ( .x(\U311/U35/Z ), .a(\U311/nz[1] ) );
    aoi222_1 \U311/U31/U30/U1  ( .x(\U311/x[1] ), .a(\net413[12] ), .b(
        \net413[13] ), .c(\net413[12] ), .d(\U311/U31/Z ), .e(\net413[13] ), 
        .f(\U311/U31/Z ) );
    inv_1 \U311/U31/U30/Uinv  ( .x(\U311/U31/Z ), .a(\U311/x[1] ) );
    aoi21_1 \U151/U30/U1/U1  ( .x(net407), .a(\U151/Z ), .b(chainff_ack), .c(
        net332) );
    inv_1 \U151/U30/U1/U2  ( .x(\U151/Z ), .a(net407) );
    ao222_1 \U324/U18/U1/U1  ( .x(hdrack), .a(ctrl_cd), .b(net383), .c(ctrl_cd
        ), .d(hdrack), .e(net383), .f(hdrack) );
    ao222_1 \U244/U18/U1/U1  ( .x(donotify), .a(done_hdr), .b(\hdr[17] ), .c(
        done_hdr), .d(donotify), .e(\hdr[17] ), .f(donotify) );
    ao222_1 \U260/U18/U1/U1  ( .x(net362), .a(net337), .b(\hdr[1] ), .c(net337
        ), .d(net362), .e(\hdr[1] ), .f(net362) );
    ao222_1 \U296/U18/U1/U1  ( .x(done_accept), .a(done_eop), .b(notify_accept
        ), .c(done_eop), .d(done_accept), .e(notify_accept), .f(done_accept)
         );
    ao222_1 \U261/U18/U1/U1  ( .x(net359), .a(net340), .b(\hdr[1] ), .c(net340
        ), .d(net359), .e(\hdr[1] ), .f(net359) );
    ao222_1 \U316/U18/U1/U1  ( .x(done_pl), .a(net364), .b(routeack), .c(
        net364), .d(done_pl), .e(routeack), .f(done_pl) );
    ao31_1 \U319/U21/U1/aoi  ( .x(\U319/U21/U1/loop ), .a(\hdr[1] ), .b(
        done_hdr), .c(rnw_h), .d(read_req) );
    oa21_1 \U319/U21/U1/outGate  ( .x(read_req), .a(\hdr[1] ), .b(done_hdr), 
        .c(\U319/U21/U1/loop ) );
    ao31_1 \U323/U21/U1/aoi  ( .x(\U323/U21/U1/loop ), .a(done_eop), .b(
        notify_defer), .c(ctrl_cd), .d(done_defer) );
    oa21_1 \U323/U21/U1/outGate  ( .x(done_defer), .a(done_eop), .b(
        notify_defer), .c(\U323/U21/U1/loop ) );
    ao31_1 \U320/U21/U1/aoi  ( .x(\U320/U21/U1/loop ), .a(\hdr[1] ), .b(
        done_hdr), .c(rnw_l), .d(dowrite) );
    oa21_1 \U320/U21/U1/outGate  ( .x(dowrite), .a(\hdr[1] ), .b(done_hdr), 
        .c(\U320/U21/U1/loop ) );
    ao31_1 \U321/U21/U1/aoi  ( .x(\U321/U21/U1/loop ), .a(read_req), .b(
        done_eop), .c(ctrl_cd), .d(done_read) );
    oa21_1 \U321/U21/U1/outGate  ( .x(done_read), .a(read_req), .b(done_eop), 
        .c(\U321/U21/U1/loop ) );
    ao31_1 \U322/U21/U1/aoi  ( .x(\U322/U21/U1/loop ), .a(dowrite), .b(
        done_eop), .c(ctrl_cd), .d(done_write) );
    oa21_1 \U322/U21/U1/outGate  ( .x(done_write), .a(dowrite), .b(done_eop), 
        .c(\U322/U21/U1/loop ) );
    nor2_2 \U210/U1703/U6  ( .x(done_hdr), .a(\U210/drivemonitor ), .b(
        \U210/naa ) );
    inv_2 \U210/U1699/U3  ( .x(\U210/net2 ), .a(\U210/net3 ) );
    and2_4 \U210/U2_0_/U8  ( .x(\drive_l[0] ), .a(net0230), .b(\U210/net2 ) );
    and2_4 \U210/U2_1_/U8  ( .x(\drive_l[1] ), .a(net0230), .b(\U210/net2 ) );
    inv_1 \U210/U1701/U3  ( .x(\U210/naa ), .a(\U210/bdone ) );
    ao222_1 \U210/U13/U18/U1/U1  ( .x(\U210/drivemonitor ), .a(\drive_l[1] ), 
        .b(\drive_l[0] ), .c(\drive_l[1] ), .d(\U210/drivemonitor ), .e(
        \drive_l[0] ), .f(\U210/drivemonitor ) );
    aoi21_1 \U210/U1702/U30/U1/U1  ( .x(\U210/bdone ), .a(\U210/U1702/Z ), .b(
        chainff_ack), .c(\U210/net2 ) );
    inv_1 \U210/U1702/U30/U1/U2  ( .x(\U210/U1702/Z ), .a(\U210/bdone ) );
    ao23_1 \U210/U1693/U21/U1/U1  ( .x(\U210/net3 ), .a(net0230), .b(
        \U210/net3 ), .c(net0230), .d(\U210/drivemonitor ), .e(chainff_ack) );
    nor2_2 \I0/U1703/U6  ( .x(net0230), .a(\I0/drivemonitor ), .b(\I0/naa ) );
    inv_2 \I0/U1699/U3  ( .x(\I0/net2 ), .a(\I0/net3 ) );
    and2_4 \I0/U2_0_/U8  ( .x(\drive_h[0] ), .a(net407), .b(\I0/net2 ) );
    and2_4 \I0/U2_1_/U8  ( .x(\drive_h[1] ), .a(net407), .b(\I0/net2 ) );
    inv_1 \I0/U1701/U3  ( .x(\I0/naa ), .a(\I0/bdone ) );
    ao222_1 \I0/U13/U18/U1/U1  ( .x(\I0/drivemonitor ), .a(\drive_h[1] ), .b(
        \drive_h[0] ), .c(\drive_h[1] ), .d(\I0/drivemonitor ), .e(
        \drive_h[0] ), .f(\I0/drivemonitor ) );
    aoi21_1 \I0/U1702/U30/U1/U1  ( .x(\I0/bdone ), .a(\I0/U1702/Z ), .b(
        chainff_ack), .c(\I0/net2 ) );
    inv_1 \I0/U1702/U30/U1/U2  ( .x(\I0/U1702/Z ), .a(\I0/bdone ) );
    ao23_1 \I0/U1693/U21/U1/U1  ( .x(\I0/net3 ), .a(net407), .b(\I0/net3 ), 
        .c(net407), .d(\I0/drivemonitor ), .e(chainff_ack) );
    buf_3 U1 ( .x(chainff_ack), .a(chainack) );
    or2_1 U2 ( .x(chainh[4]), .a(chain_ff_h[4]), .b(\net284[3] ) );
    or2_1 U3 ( .x(chainh[2]), .a(chain_ff_h[2]), .b(\net284[5] ) );
    or2_1 U4 ( .x(chainl[3]), .a(chainff_l[3]), .b(\net288[4] ) );
endmodule


module chain_tchdr_2 ( addr_req, col_h, col_l, itag_h, itag_l, lock, ncback, 
    neop, pred, pullcd, reset, rnw_h, rnw_l, seq, size_h, size_l, write_req, 
    chwh, chwl, addr_ack, addr_pull, nReset, nack, write_ack, write_pull );
output [2:0] col_h;
output [2:0] col_l;
output [4:0] itag_h;
output [4:0] itag_l;
output [1:0] lock;
output [1:0] pred;
output [1:0] seq;
output [1:0] size_h;
output [1:0] size_l;
input  [7:0] chwh;
input  [7:0] chwl;
input  addr_ack, addr_pull, nReset, nack, write_ack, write_pull;
output addr_req, ncback, neop, pullcd, reset, rnw_h, rnw_l, write_req;
    wire \ncd[7] , \ncd[6] , \ncd[5] , \ncd[4] , \ncd[3] , \ncd[2] , \ncd[1] , 
        \ncd[0] , net88, receive, pullcdwk, read, net83, ack, net94, n9, 
        \U1664/U28/Z , \U1664/U32/Z , \U1664/U29/Z , \U1664/U33/Z , 
        \U1664/U30/Z , \U1664/U31/Z , \U1664/U37/Z , \U473/Z , \U1664/y[0] , 
        \U1664/y[1] , \U1664/x[1] , \U1664/x[3] , \U1664/x[2] , \U1664/x[0] , 
        \hdr_hld/oh[4] , \hdr_hld/oh[3] , \hdr_hld/ol[4] , \hdr_hld/ol[3] , 
        \hdr_hld/net20 , \hdr_hld/net33 , \hdr_hld/net32 , 
        \hdr_hld/low/drivel , \hdr_hld/low/driveh , \hdr_hld/low/localcd , 
        \hdr_hld/low/ncd[7] , \hdr_hld/low/ncd[6] , \hdr_hld/low/ncd[5] , 
        \hdr_hld/low/ncd[4] , \hdr_hld/low/ncd[3] , \hdr_hld/low/ncd[2] , 
        \hdr_hld/low/ncd[1] , \hdr_hld/low/ncd[0] , \hdr_hld/low/ba , 
        \hdr_hld/low/latch , \hdr_hld/low/acb , \hdr_hld/low/ctrlack_internal , 
        \hdr_hld/low/nlocalcd , \hdr_hld/low/U4/U28/U1/clr , 
        \hdr_hld/low/U4/U28/U1/set , \hdr_hld/low/U1/Z , 
        \hdr_hld/low/U1664/y[0] , \hdr_hld/low/U1664/y[1] , 
        \hdr_hld/low/U1664/x[1] , \hdr_hld/low/U1664/x[3] , 
        \hdr_hld/low/U1664/x[2] , \hdr_hld/low/U1664/x[0] , 
        \hdr_hld/low/U1664/U28/Z , \hdr_hld/low/U1664/U32/Z , 
        \hdr_hld/low/U1664/U29/Z , \hdr_hld/low/U1664/U33/Z , 
        \hdr_hld/low/U1664/U30/Z , \hdr_hld/low/U1664/U31/Z , 
        \hdr_hld/low/U1664/U37/Z , \hdr_hld/low/U1669/nr , 
        \hdr_hld/low/U1669/nd , \hdr_hld/low/U1669/n2 , \hdr_hld/high/drivel , 
        \hdr_hld/high/driveh , \hdr_hld/high/localcd , \hdr_hld/high/ncd[7] , 
        \hdr_hld/high/ncd[6] , \hdr_hld/high/ncd[5] , \hdr_hld/high/ncd[4] , 
        \hdr_hld/high/ncd[3] , \hdr_hld/high/ncd[2] , \hdr_hld/high/ncd[1] , 
        \hdr_hld/high/ncd[0] , \hdr_hld/high/ba , \hdr_hld/high/latch , 
        \hdr_hld/high/acb , \hdr_hld/high/ctrlack_internal , 
        \hdr_hld/high/nlocalcd , \hdr_hld/high/U4/U28/U1/clr , 
        \hdr_hld/high/U4/U28/U1/set , \hdr_hld/high/U1/Z , 
        \hdr_hld/high/U1664/y[0] , \hdr_hld/high/U1664/y[1] , 
        \hdr_hld/high/U1664/x[1] , \hdr_hld/high/U1664/x[3] , 
        \hdr_hld/high/U1664/x[2] , \hdr_hld/high/U1664/x[0] , 
        \hdr_hld/high/U1664/U28/Z , \hdr_hld/high/U1664/U32/Z , 
        \hdr_hld/high/U1664/U29/Z , \hdr_hld/high/U1664/U33/Z , 
        \hdr_hld/high/U1664/U30/Z , \hdr_hld/high/U1664/U31/Z , 
        \hdr_hld/high/U1664/U37/Z , \hdr_hld/high/U1669/nr , 
        \hdr_hld/high/U1669/nd , \hdr_hld/high/U1669/n2 , n1, n2, n3, n4, n5, 
        n6, n7;
    buf_1 U262 ( .x(n9), .a(pullcdwk) );
    or3_2 \U1668/U12  ( .x(ncback), .a(net94), .b(addr_pull), .c(write_pull)
         );
    inv_1 \I0/U3  ( .x(net94), .a(net88) );
    nor2_1 \U514_0_/U5  ( .x(\ncd[0] ), .a(chwh[0]), .b(chwl[0]) );
    nor2_1 \U514_1_/U5  ( .x(\ncd[1] ), .a(chwh[1]), .b(chwl[1]) );
    nor2_1 \U514_2_/U5  ( .x(\ncd[2] ), .a(chwh[2]), .b(chwl[2]) );
    nor2_1 \U514_3_/U5  ( .x(\ncd[3] ), .a(chwh[3]), .b(chwl[3]) );
    nor2_1 \U514_4_/U5  ( .x(\ncd[4] ), .a(chwh[4]), .b(chwl[4]) );
    nor2_1 \U514_5_/U5  ( .x(\ncd[5] ), .a(chwh[5]), .b(chwl[5]) );
    nor2_1 \U514_6_/U5  ( .x(\ncd[6] ), .a(chwh[6]), .b(chwl[6]) );
    nor2_1 \U514_7_/U5  ( .x(\ncd[7] ), .a(chwh[7]), .b(chwl[7]) );
    nor2_1 \U1669/U5  ( .x(neop), .a(read), .b(write_ack) );
    nand2_1 \U303/U5  ( .x(ack), .a(nack), .b(nReset) );
    nand2_1 \U1670/U5  ( .x(net83), .a(neop), .b(nReset) );
    ao222_1 \U47/U18/U1/U1  ( .x(read), .a(addr_ack), .b(rnw_h), .c(addr_ack), 
        .d(read), .e(rnw_h), .f(read) );
    ao222_1 \U48/U18/U1/U1  ( .x(write_req), .a(rnw_l), .b(addr_ack), .c(rnw_l
        ), .d(write_req), .e(addr_ack), .f(write_req) );
    aoi222_1 \U1664/U28/U30/U1  ( .x(\U1664/x[3] ), .a(\ncd[7] ), .b(\ncd[6] ), 
        .c(\ncd[7] ), .d(\U1664/U28/Z ), .e(\ncd[6] ), .f(\U1664/U28/Z ) );
    inv_1 \U1664/U28/U30/Uinv  ( .x(\U1664/U28/Z ), .a(\U1664/x[3] ) );
    aoi222_1 \U1664/U32/U30/U1  ( .x(\U1664/x[0] ), .a(\ncd[1] ), .b(\ncd[0] ), 
        .c(\ncd[1] ), .d(\U1664/U32/Z ), .e(\ncd[0] ), .f(\U1664/U32/Z ) );
    inv_1 \U1664/U32/U30/Uinv  ( .x(\U1664/U32/Z ), .a(\U1664/x[0] ) );
    aoi222_1 \U1664/U29/U30/U1  ( .x(\U1664/x[2] ), .a(\ncd[5] ), .b(\ncd[4] ), 
        .c(\ncd[5] ), .d(\U1664/U29/Z ), .e(\ncd[4] ), .f(\U1664/U29/Z ) );
    inv_1 \U1664/U29/U30/Uinv  ( .x(\U1664/U29/Z ), .a(\U1664/x[2] ) );
    aoi222_1 \U1664/U33/U30/U1  ( .x(\U1664/y[0] ), .a(\U1664/x[1] ), .b(
        \U1664/x[0] ), .c(\U1664/x[1] ), .d(\U1664/U33/Z ), .e(\U1664/x[0] ), 
        .f(\U1664/U33/Z ) );
    inv_1 \U1664/U33/U30/Uinv  ( .x(\U1664/U33/Z ), .a(\U1664/y[0] ) );
    aoi222_1 \U1664/U30/U30/U1  ( .x(\U1664/y[1] ), .a(\U1664/x[3] ), .b(
        \U1664/x[2] ), .c(\U1664/x[3] ), .d(\U1664/U30/Z ), .e(\U1664/x[2] ), 
        .f(\U1664/U30/Z ) );
    inv_1 \U1664/U30/U30/Uinv  ( .x(\U1664/U30/Z ), .a(\U1664/y[1] ) );
    aoi222_1 \U1664/U31/U30/U1  ( .x(\U1664/x[1] ), .a(\ncd[3] ), .b(\ncd[2] ), 
        .c(\ncd[3] ), .d(\U1664/U31/Z ), .e(\ncd[2] ), .f(\U1664/U31/Z ) );
    inv_1 \U1664/U31/U30/Uinv  ( .x(\U1664/U31/Z ), .a(\U1664/x[1] ) );
    aoi222_1 \U1664/U37/U30/U1  ( .x(pullcdwk), .a(\U1664/y[0] ), .b(
        \U1664/y[1] ), .c(\U1664/y[0] ), .d(\U1664/U37/Z ), .e(\U1664/y[1] ), 
        .f(\U1664/U37/Z ) );
    inv_1 \U1664/U37/U30/Uinv  ( .x(\U1664/U37/Z ), .a(pullcdwk) );
    aoi222_1 \U473/U30/U1  ( .x(receive), .a(net83), .b(ack), .c(net83), .d(
        \U473/Z ), .e(ack), .f(\U473/Z ) );
    inv_1 \U473/U30/Uinv  ( .x(\U473/Z ), .a(receive) );
    nor2_1 \hdr_hld/U3/U5  ( .x(net88), .a(\hdr_hld/net32 ), .b(
        \hdr_hld/net33 ) );
    buf_2 \hdr_hld/low/U1653  ( .x(\hdr_hld/low/latch ), .a(\hdr_hld/net32 )
         );
    nor2_1 \hdr_hld/low/U264/U5  ( .x(\hdr_hld/low/nlocalcd ), .a(reset), .b(
        \hdr_hld/low/localcd ) );
    nor2_1 \hdr_hld/low/U1659_0_/U5  ( .x(\hdr_hld/low/ncd[0] ), .a(seq[0]), 
        .b(seq[1]) );
    nor2_1 \hdr_hld/low/U1659_1_/U5  ( .x(\hdr_hld/low/ncd[1] ), .a(pred[0]), 
        .b(pred[1]) );
    nor2_1 \hdr_hld/low/U1659_2_/U5  ( .x(\hdr_hld/low/ncd[2] ), .a(lock[0]), 
        .b(lock[1]) );
    nor2_1 \hdr_hld/low/U1659_3_/U5  ( .x(\hdr_hld/low/ncd[3] ), .a(
        \hdr_hld/ol[3] ), .b(\hdr_hld/oh[3] ) );
    nor2_1 \hdr_hld/low/U1659_4_/U5  ( .x(\hdr_hld/low/ncd[4] ), .a(
        \hdr_hld/ol[4] ), .b(\hdr_hld/oh[4] ) );
    nor2_1 \hdr_hld/low/U1659_5_/U5  ( .x(\hdr_hld/low/ncd[5] ), .a(rnw_l), 
        .b(rnw_h) );
    nor2_1 \hdr_hld/low/U1659_6_/U5  ( .x(\hdr_hld/low/ncd[6] ), .a(size_l[0]), 
        .b(size_h[0]) );
    nor2_1 \hdr_hld/low/U1659_7_/U5  ( .x(\hdr_hld/low/ncd[7] ), .a(size_l[1]), 
        .b(size_h[1]) );
    nor2_1 \hdr_hld/low/U3/U5  ( .x(\hdr_hld/low/ctrlack_internal ), .a(
        \hdr_hld/low/acb ), .b(\hdr_hld/low/ba ) );
    buf_2 \hdr_hld/low/U1665/U7  ( .x(\hdr_hld/low/driveh ), .a(
        \hdr_hld/net20 ) );
    buf_2 \hdr_hld/low/U1666/U7  ( .x(\hdr_hld/low/drivel ), .a(
        \hdr_hld/net20 ) );
    ao23_1 \hdr_hld/low/U1658_0_/U21/U1/U1  ( .x(seq[0]), .a(n2), .b(seq[0]), 
        .c(\hdr_hld/low/drivel ), .d(chwl[0]), .e(n3) );
    ao23_1 \hdr_hld/low/U1658_1_/U21/U1/U1  ( .x(pred[0]), .a(n1), .b(pred[0]), 
        .c(\hdr_hld/low/drivel ), .d(chwl[1]), .e(n3) );
    ao23_1 \hdr_hld/low/U1658_2_/U21/U1/U1  ( .x(lock[0]), .a(n1), .b(lock[0]), 
        .c(\hdr_hld/low/driveh ), .d(chwl[2]), .e(n3) );
    ao23_1 \hdr_hld/low/U1658_3_/U21/U1/U1  ( .x(\hdr_hld/ol[3] ), .a(n1), .b(
        \hdr_hld/ol[3] ), .c(\hdr_hld/low/driveh ), .d(chwl[3]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_4_/U21/U1/U1  ( .x(\hdr_hld/ol[4] ), .a(n2), .b(
        \hdr_hld/ol[4] ), .c(\hdr_hld/low/drivel ), .d(chwl[4]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_5_/U21/U1/U1  ( .x(rnw_l), .a(
        \hdr_hld/low/driveh ), .b(rnw_l), .c(\hdr_hld/low/driveh ), .d(chwl[5]
        ), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_6_/U21/U1/U1  ( .x(size_l[0]), .a(
        \hdr_hld/low/drivel ), .b(size_l[0]), .c(n2), .d(chwl[6]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_7_/U21/U1/U1  ( .x(size_l[1]), .a(
        \hdr_hld/low/drivel ), .b(size_l[1]), .c(\hdr_hld/low/drivel ), .d(
        chwl[7]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_0_/U21/U1/U1  ( .x(seq[1]), .a(
        \hdr_hld/low/drivel ), .b(seq[1]), .c(\hdr_hld/low/driveh ), .d(chwh
        [0]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_1_/U21/U1/U1  ( .x(pred[1]), .a(
        \hdr_hld/low/driveh ), .b(pred[1]), .c(n1), .d(chwh[1]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_2_/U21/U1/U1  ( .x(lock[1]), .a(
        \hdr_hld/low/driveh ), .b(lock[1]), .c(n1), .d(chwh[2]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_3_/U21/U1/U1  ( .x(\hdr_hld/oh[3] ), .a(
        \hdr_hld/low/drivel ), .b(\hdr_hld/oh[3] ), .c(n2), .d(chwh[3]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_4_/U21/U1/U1  ( .x(\hdr_hld/oh[4] ), .a(n2), .b(
        \hdr_hld/oh[4] ), .c(n1), .d(chwh[4]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_5_/U21/U1/U1  ( .x(rnw_h), .a(n2), .b(rnw_h), 
        .c(n1), .d(chwh[5]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_6_/U21/U1/U1  ( .x(size_h[0]), .a(n1), .b(size_h
        [0]), .c(n2), .d(chwh[6]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_7_/U21/U1/U1  ( .x(size_h[1]), .a(
        \hdr_hld/low/driveh ), .b(size_h[1]), .c(n2), .d(chwh[7]), .e(
        \hdr_hld/low/latch ) );
    aoai211_1 \hdr_hld/low/U4/U28/U1/U1  ( .x(\hdr_hld/low/U4/U28/U1/clr ), 
        .a(\hdr_hld/net20 ), .b(\hdr_hld/low/acb ), .c(\hdr_hld/low/nlocalcd ), 
        .d(\hdr_hld/net32 ) );
    nand3_1 \hdr_hld/low/U4/U28/U1/U2  ( .x(\hdr_hld/low/U4/U28/U1/set ), .a(
        \hdr_hld/low/nlocalcd ), .b(\hdr_hld/net20 ), .c(\hdr_hld/low/acb ) );
    nand2_2 \hdr_hld/low/U4/U28/U1/U3  ( .x(\hdr_hld/net32 ), .a(
        \hdr_hld/low/U4/U28/U1/clr ), .b(\hdr_hld/low/U4/U28/U1/set ) );
    oai21_1 \hdr_hld/low/U1/U30/U1/U1  ( .x(\hdr_hld/low/acb ), .a(
        \hdr_hld/low/U1/Z ), .b(\hdr_hld/low/ba ), .c(\hdr_hld/net20 ) );
    inv_1 \hdr_hld/low/U1/U30/U1/U2  ( .x(\hdr_hld/low/U1/Z ), .a(
        \hdr_hld/low/acb ) );
    ao222_1 \hdr_hld/low/U5/U18/U1/U1  ( .x(\hdr_hld/low/ba ), .a(
        \hdr_hld/low/latch ), .b(n9), .c(\hdr_hld/low/latch ), .d(
        \hdr_hld/low/ba ), .e(n9), .f(\hdr_hld/low/ba ) );
    aoi222_1 \hdr_hld/low/U1664/U28/U30/U1  ( .x(\hdr_hld/low/U1664/x[3] ), 
        .a(\hdr_hld/low/ncd[7] ), .b(\hdr_hld/low/ncd[6] ), .c(
        \hdr_hld/low/ncd[7] ), .d(\hdr_hld/low/U1664/U28/Z ), .e(
        \hdr_hld/low/ncd[6] ), .f(\hdr_hld/low/U1664/U28/Z ) );
    inv_1 \hdr_hld/low/U1664/U28/U30/Uinv  ( .x(\hdr_hld/low/U1664/U28/Z ), 
        .a(\hdr_hld/low/U1664/x[3] ) );
    aoi222_1 \hdr_hld/low/U1664/U32/U30/U1  ( .x(\hdr_hld/low/U1664/x[0] ), 
        .a(\hdr_hld/low/ncd[1] ), .b(\hdr_hld/low/ncd[0] ), .c(
        \hdr_hld/low/ncd[1] ), .d(\hdr_hld/low/U1664/U32/Z ), .e(
        \hdr_hld/low/ncd[0] ), .f(\hdr_hld/low/U1664/U32/Z ) );
    inv_1 \hdr_hld/low/U1664/U32/U30/Uinv  ( .x(\hdr_hld/low/U1664/U32/Z ), 
        .a(\hdr_hld/low/U1664/x[0] ) );
    aoi222_1 \hdr_hld/low/U1664/U29/U30/U1  ( .x(\hdr_hld/low/U1664/x[2] ), 
        .a(\hdr_hld/low/ncd[5] ), .b(\hdr_hld/low/ncd[4] ), .c(
        \hdr_hld/low/ncd[5] ), .d(\hdr_hld/low/U1664/U29/Z ), .e(
        \hdr_hld/low/ncd[4] ), .f(\hdr_hld/low/U1664/U29/Z ) );
    inv_1 \hdr_hld/low/U1664/U29/U30/Uinv  ( .x(\hdr_hld/low/U1664/U29/Z ), 
        .a(\hdr_hld/low/U1664/x[2] ) );
    aoi222_1 \hdr_hld/low/U1664/U33/U30/U1  ( .x(\hdr_hld/low/U1664/y[0] ), 
        .a(\hdr_hld/low/U1664/x[1] ), .b(\hdr_hld/low/U1664/x[0] ), .c(
        \hdr_hld/low/U1664/x[1] ), .d(\hdr_hld/low/U1664/U33/Z ), .e(
        \hdr_hld/low/U1664/x[0] ), .f(\hdr_hld/low/U1664/U33/Z ) );
    inv_1 \hdr_hld/low/U1664/U33/U30/Uinv  ( .x(\hdr_hld/low/U1664/U33/Z ), 
        .a(\hdr_hld/low/U1664/y[0] ) );
    aoi222_1 \hdr_hld/low/U1664/U30/U30/U1  ( .x(\hdr_hld/low/U1664/y[1] ), 
        .a(\hdr_hld/low/U1664/x[3] ), .b(\hdr_hld/low/U1664/x[2] ), .c(
        \hdr_hld/low/U1664/x[3] ), .d(\hdr_hld/low/U1664/U30/Z ), .e(
        \hdr_hld/low/U1664/x[2] ), .f(\hdr_hld/low/U1664/U30/Z ) );
    inv_1 \hdr_hld/low/U1664/U30/U30/Uinv  ( .x(\hdr_hld/low/U1664/U30/Z ), 
        .a(\hdr_hld/low/U1664/y[1] ) );
    aoi222_1 \hdr_hld/low/U1664/U31/U30/U1  ( .x(\hdr_hld/low/U1664/x[1] ), 
        .a(\hdr_hld/low/ncd[3] ), .b(\hdr_hld/low/ncd[2] ), .c(
        \hdr_hld/low/ncd[3] ), .d(\hdr_hld/low/U1664/U31/Z ), .e(
        \hdr_hld/low/ncd[2] ), .f(\hdr_hld/low/U1664/U31/Z ) );
    inv_1 \hdr_hld/low/U1664/U31/U30/Uinv  ( .x(\hdr_hld/low/U1664/U31/Z ), 
        .a(\hdr_hld/low/U1664/x[1] ) );
    aoi222_1 \hdr_hld/low/U1664/U37/U30/U1  ( .x(\hdr_hld/low/localcd ), .a(
        \hdr_hld/low/U1664/y[0] ), .b(\hdr_hld/low/U1664/y[1] ), .c(
        \hdr_hld/low/U1664/y[0] ), .d(\hdr_hld/low/U1664/U37/Z ), .e(
        \hdr_hld/low/U1664/y[1] ), .f(\hdr_hld/low/U1664/U37/Z ) );
    inv_1 \hdr_hld/low/U1664/U37/U30/Uinv  ( .x(\hdr_hld/low/U1664/U37/Z ), 
        .a(\hdr_hld/low/localcd ) );
    nor3_1 \hdr_hld/low/U1669/Unr  ( .x(\hdr_hld/low/U1669/nr ), .a(
        \hdr_hld/low/ctrlack_internal ), .b(\hdr_hld/low/driveh ), .c(n1) );
    nand3_1 \hdr_hld/low/U1669/Und  ( .x(\hdr_hld/low/U1669/nd ), .a(
        \hdr_hld/low/ctrlack_internal ), .b(n2), .c(\hdr_hld/low/drivel ) );
    oa21_1 \hdr_hld/low/U1669/U1  ( .x(\hdr_hld/low/U1669/n2 ), .a(
        \hdr_hld/low/U1669/n2 ), .b(\hdr_hld/low/U1669/nr ), .c(
        \hdr_hld/low/U1669/nd ) );
    inv_2 \hdr_hld/low/U1669/U3  ( .x(addr_req), .a(\hdr_hld/low/U1669/n2 ) );
    buf_2 \hdr_hld/high/U1653  ( .x(\hdr_hld/high/latch ), .a(\hdr_hld/net33 )
         );
    nor2_1 \hdr_hld/high/U264/U5  ( .x(\hdr_hld/high/nlocalcd ), .a(reset), 
        .b(\hdr_hld/high/localcd ) );
    nor2_1 \hdr_hld/high/U1659_0_/U5  ( .x(\hdr_hld/high/ncd[0] ), .a(itag_l
        [0]), .b(itag_h[0]) );
    nor2_1 \hdr_hld/high/U1659_1_/U5  ( .x(\hdr_hld/high/ncd[1] ), .a(itag_l
        [1]), .b(itag_h[1]) );
    nor2_1 \hdr_hld/high/U1659_2_/U5  ( .x(\hdr_hld/high/ncd[2] ), .a(itag_l
        [2]), .b(itag_h[2]) );
    nor2_1 \hdr_hld/high/U1659_3_/U5  ( .x(\hdr_hld/high/ncd[3] ), .a(itag_l
        [3]), .b(itag_h[3]) );
    nor2_1 \hdr_hld/high/U1659_4_/U5  ( .x(\hdr_hld/high/ncd[4] ), .a(itag_l
        [4]), .b(itag_h[4]) );
    nor2_1 \hdr_hld/high/U1659_5_/U5  ( .x(\hdr_hld/high/ncd[5] ), .a(col_l[0]
        ), .b(col_h[0]) );
    nor2_1 \hdr_hld/high/U1659_6_/U5  ( .x(\hdr_hld/high/ncd[6] ), .a(col_l[1]
        ), .b(col_h[1]) );
    nor2_1 \hdr_hld/high/U1659_7_/U5  ( .x(\hdr_hld/high/ncd[7] ), .a(col_l[2]
        ), .b(col_h[2]) );
    nor2_1 \hdr_hld/high/U3/U5  ( .x(\hdr_hld/high/ctrlack_internal ), .a(
        \hdr_hld/high/acb ), .b(\hdr_hld/high/ba ) );
    buf_2 \hdr_hld/high/U1665/U7  ( .x(\hdr_hld/high/driveh ), .a(receive) );
    buf_2 \hdr_hld/high/U1666/U7  ( .x(\hdr_hld/high/drivel ), .a(receive) );
    ao23_1 \hdr_hld/high/U1658_0_/U21/U1/U1  ( .x(itag_l[0]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[0]), .c(\hdr_hld/high/drivel ), .d(
        chwl[0]), .e(n7) );
    ao23_1 \hdr_hld/high/U1658_1_/U21/U1/U1  ( .x(itag_l[1]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[1]), .c(\hdr_hld/high/drivel ), .d(
        chwl[1]), .e(n7) );
    ao23_1 \hdr_hld/high/U1658_2_/U21/U1/U1  ( .x(itag_l[2]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[2]), .c(\hdr_hld/high/drivel ), .d(
        chwl[2]), .e(n7) );
    ao23_1 \hdr_hld/high/U1658_3_/U21/U1/U1  ( .x(itag_l[3]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[3]), .c(\hdr_hld/high/drivel ), .d(
        chwl[3]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1658_4_/U21/U1/U1  ( .x(itag_l[4]), .a(n4), .b(
        itag_l[4]), .c(\hdr_hld/high/drivel ), .d(chwl[4]), .e(
        \hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1658_5_/U21/U1/U1  ( .x(col_l[0]), .a(n4), .b(col_l
        [0]), .c(\hdr_hld/high/drivel ), .d(chwl[5]), .e(\hdr_hld/high/latch )
         );
    ao23_1 \hdr_hld/high/U1658_6_/U21/U1/U1  ( .x(col_l[1]), .a(
        \hdr_hld/high/drivel ), .b(col_l[1]), .c(\hdr_hld/high/drivel ), .d(
        chwl[6]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1658_7_/U21/U1/U1  ( .x(col_l[2]), .a(n4), .b(col_l
        [2]), .c(\hdr_hld/high/drivel ), .d(chwl[7]), .e(\hdr_hld/high/latch )
         );
    ao23_1 \hdr_hld/high/U1651_0_/U21/U1/U1  ( .x(itag_h[0]), .a(n5), .b(
        itag_h[0]), .c(n5), .d(chwh[0]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_1_/U21/U1/U1  ( .x(itag_h[1]), .a(n5), .b(
        itag_h[1]), .c(n6), .d(chwh[1]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_2_/U21/U1/U1  ( .x(itag_h[2]), .a(n5), .b(
        itag_h[2]), .c(n6), .d(chwh[2]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_3_/U21/U1/U1  ( .x(itag_h[3]), .a(n5), .b(
        itag_h[3]), .c(n6), .d(chwh[3]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_4_/U21/U1/U1  ( .x(itag_h[4]), .a(n5), .b(
        itag_h[4]), .c(n6), .d(chwh[4]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_5_/U21/U1/U1  ( .x(col_h[0]), .a(n5), .b(col_h
        [0]), .c(n6), .d(chwh[5]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_6_/U21/U1/U1  ( .x(col_h[1]), .a(n5), .b(col_h
        [1]), .c(n5), .d(chwh[6]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_7_/U21/U1/U1  ( .x(col_h[2]), .a(n5), .b(col_h
        [2]), .c(n5), .d(chwh[7]), .e(\hdr_hld/high/latch ) );
    aoai211_1 \hdr_hld/high/U4/U28/U1/U1  ( .x(\hdr_hld/high/U4/U28/U1/clr ), 
        .a(receive), .b(\hdr_hld/high/acb ), .c(\hdr_hld/high/nlocalcd ), .d(
        \hdr_hld/net33 ) );
    nand3_1 \hdr_hld/high/U4/U28/U1/U2  ( .x(\hdr_hld/high/U4/U28/U1/set ), 
        .a(\hdr_hld/high/nlocalcd ), .b(receive), .c(\hdr_hld/high/acb ) );
    nand2_2 \hdr_hld/high/U4/U28/U1/U3  ( .x(\hdr_hld/net33 ), .a(
        \hdr_hld/high/U4/U28/U1/clr ), .b(\hdr_hld/high/U4/U28/U1/set ) );
    oai21_1 \hdr_hld/high/U1/U30/U1/U1  ( .x(\hdr_hld/high/acb ), .a(
        \hdr_hld/high/U1/Z ), .b(\hdr_hld/high/ba ), .c(receive) );
    inv_1 \hdr_hld/high/U1/U30/U1/U2  ( .x(\hdr_hld/high/U1/Z ), .a(
        \hdr_hld/high/acb ) );
    ao222_1 \hdr_hld/high/U5/U18/U1/U1  ( .x(\hdr_hld/high/ba ), .a(
        \hdr_hld/high/latch ), .b(n9), .c(\hdr_hld/high/latch ), .d(
        \hdr_hld/high/ba ), .e(n9), .f(\hdr_hld/high/ba ) );
    aoi222_1 \hdr_hld/high/U1664/U28/U30/U1  ( .x(\hdr_hld/high/U1664/x[3] ), 
        .a(\hdr_hld/high/ncd[7] ), .b(\hdr_hld/high/ncd[6] ), .c(
        \hdr_hld/high/ncd[7] ), .d(\hdr_hld/high/U1664/U28/Z ), .e(
        \hdr_hld/high/ncd[6] ), .f(\hdr_hld/high/U1664/U28/Z ) );
    inv_1 \hdr_hld/high/U1664/U28/U30/Uinv  ( .x(\hdr_hld/high/U1664/U28/Z ), 
        .a(\hdr_hld/high/U1664/x[3] ) );
    aoi222_1 \hdr_hld/high/U1664/U32/U30/U1  ( .x(\hdr_hld/high/U1664/x[0] ), 
        .a(\hdr_hld/high/ncd[1] ), .b(\hdr_hld/high/ncd[0] ), .c(
        \hdr_hld/high/ncd[1] ), .d(\hdr_hld/high/U1664/U32/Z ), .e(
        \hdr_hld/high/ncd[0] ), .f(\hdr_hld/high/U1664/U32/Z ) );
    inv_1 \hdr_hld/high/U1664/U32/U30/Uinv  ( .x(\hdr_hld/high/U1664/U32/Z ), 
        .a(\hdr_hld/high/U1664/x[0] ) );
    aoi222_1 \hdr_hld/high/U1664/U29/U30/U1  ( .x(\hdr_hld/high/U1664/x[2] ), 
        .a(\hdr_hld/high/ncd[5] ), .b(\hdr_hld/high/ncd[4] ), .c(
        \hdr_hld/high/ncd[5] ), .d(\hdr_hld/high/U1664/U29/Z ), .e(
        \hdr_hld/high/ncd[4] ), .f(\hdr_hld/high/U1664/U29/Z ) );
    inv_1 \hdr_hld/high/U1664/U29/U30/Uinv  ( .x(\hdr_hld/high/U1664/U29/Z ), 
        .a(\hdr_hld/high/U1664/x[2] ) );
    aoi222_1 \hdr_hld/high/U1664/U33/U30/U1  ( .x(\hdr_hld/high/U1664/y[0] ), 
        .a(\hdr_hld/high/U1664/x[1] ), .b(\hdr_hld/high/U1664/x[0] ), .c(
        \hdr_hld/high/U1664/x[1] ), .d(\hdr_hld/high/U1664/U33/Z ), .e(
        \hdr_hld/high/U1664/x[0] ), .f(\hdr_hld/high/U1664/U33/Z ) );
    inv_1 \hdr_hld/high/U1664/U33/U30/Uinv  ( .x(\hdr_hld/high/U1664/U33/Z ), 
        .a(\hdr_hld/high/U1664/y[0] ) );
    aoi222_1 \hdr_hld/high/U1664/U30/U30/U1  ( .x(\hdr_hld/high/U1664/y[1] ), 
        .a(\hdr_hld/high/U1664/x[3] ), .b(\hdr_hld/high/U1664/x[2] ), .c(
        \hdr_hld/high/U1664/x[3] ), .d(\hdr_hld/high/U1664/U30/Z ), .e(
        \hdr_hld/high/U1664/x[2] ), .f(\hdr_hld/high/U1664/U30/Z ) );
    inv_1 \hdr_hld/high/U1664/U30/U30/Uinv  ( .x(\hdr_hld/high/U1664/U30/Z ), 
        .a(\hdr_hld/high/U1664/y[1] ) );
    aoi222_1 \hdr_hld/high/U1664/U31/U30/U1  ( .x(\hdr_hld/high/U1664/x[1] ), 
        .a(\hdr_hld/high/ncd[3] ), .b(\hdr_hld/high/ncd[2] ), .c(
        \hdr_hld/high/ncd[3] ), .d(\hdr_hld/high/U1664/U31/Z ), .e(
        \hdr_hld/high/ncd[2] ), .f(\hdr_hld/high/U1664/U31/Z ) );
    inv_1 \hdr_hld/high/U1664/U31/U30/Uinv  ( .x(\hdr_hld/high/U1664/U31/Z ), 
        .a(\hdr_hld/high/U1664/x[1] ) );
    aoi222_1 \hdr_hld/high/U1664/U37/U30/U1  ( .x(\hdr_hld/high/localcd ), .a(
        \hdr_hld/high/U1664/y[0] ), .b(\hdr_hld/high/U1664/y[1] ), .c(
        \hdr_hld/high/U1664/y[0] ), .d(\hdr_hld/high/U1664/U37/Z ), .e(
        \hdr_hld/high/U1664/y[1] ), .f(\hdr_hld/high/U1664/U37/Z ) );
    inv_1 \hdr_hld/high/U1664/U37/U30/Uinv  ( .x(\hdr_hld/high/U1664/U37/Z ), 
        .a(\hdr_hld/high/localcd ) );
    nor3_1 \hdr_hld/high/U1669/Unr  ( .x(\hdr_hld/high/U1669/nr ), .a(
        \hdr_hld/high/ctrlack_internal ), .b(\hdr_hld/high/drivel ), .c(n6) );
    nand3_1 \hdr_hld/high/U1669/Und  ( .x(\hdr_hld/high/U1669/nd ), .a(
        \hdr_hld/high/ctrlack_internal ), .b(\hdr_hld/high/drivel ), .c(n6) );
    oa21_1 \hdr_hld/high/U1669/U1  ( .x(\hdr_hld/high/U1669/n2 ), .a(
        \hdr_hld/high/U1669/n2 ), .b(\hdr_hld/high/U1669/nr ), .c(
        \hdr_hld/high/U1669/nd ) );
    inv_2 \hdr_hld/high/U1669/U3  ( .x(\hdr_hld/net20 ), .a(
        \hdr_hld/high/U1669/n2 ) );
    buf_2 U1 ( .x(n2), .a(\hdr_hld/net20 ) );
    buf_2 U2 ( .x(n1), .a(\hdr_hld/net20 ) );
    buf_1 U3 ( .x(n3), .a(\hdr_hld/low/latch ) );
    buf_1 U4 ( .x(n4), .a(\hdr_hld/high/drivel ) );
    buf_3 U5 ( .x(n5), .a(\hdr_hld/high/driveh ) );
    buf_3 U6 ( .x(n6), .a(\hdr_hld/high/driveh ) );
    buf_1 U7 ( .x(n7), .a(\hdr_hld/high/latch ) );
    inv_2 U8 ( .x(reset), .a(nReset) );
    buf_3 U9 ( .x(pullcd), .a(n9) );
endmodule


module chain_irdemux_32new_4 ( ctrlack, oh, ol, pullreq, pull_h, pull_l, 
    pullcd, reset, ctrlreq );
output [31:0] oh;
output [31:0] ol;
input  [7:0] pull_h;
input  [7:0] pull_l;
input  pullcd, reset, ctrlreq;
output ctrlack, pullreq;
    wire net30, net31, net17, \I0/net20 , \I0/net33 , \I0/net32 , 
        \I0/low/drivel , \I0/low/driveh , \I0/low/localcd , \I0/low/ncd[7] , 
        \I0/low/ncd[6] , \I0/low/ncd[5] , \I0/low/ncd[4] , \I0/low/ncd[3] , 
        \I0/low/ncd[2] , \I0/low/ncd[1] , \I0/low/ncd[0] , \I0/low/ba , 
        \I0/low/latch , \I0/low/acb , \I0/low/ctrlack_internal , 
        \I0/low/nlocalcd , \I0/low/U4/U28/U1/clr , \I0/low/U4/U28/U1/set , 
        \I0/low/U1/Z , \I0/low/U1664/y[0] , \I0/low/U1664/y[1] , 
        \I0/low/U1664/x[1] , \I0/low/U1664/x[3] , \I0/low/U1664/x[2] , 
        \I0/low/U1664/x[0] , \I0/low/U1664/U28/Z , \I0/low/U1664/U32/Z , 
        \I0/low/U1664/U29/Z , \I0/low/U1664/U33/Z , \I0/low/U1664/U30/Z , 
        \I0/low/U1664/U31/Z , \I0/low/U1664/U37/Z , \I0/low/U1669/nr , 
        \I0/low/U1669/nd , \I0/low/U1669/n2 , \I0/high/drivel , 
        \I0/high/driveh , \I0/high/localcd , \I0/high/ncd[7] , 
        \I0/high/ncd[6] , \I0/high/ncd[5] , \I0/high/ncd[4] , \I0/high/ncd[3] , 
        \I0/high/ncd[2] , \I0/high/ncd[1] , \I0/high/ncd[0] , \I0/high/ba , 
        \I0/high/latch , \I0/high/acb , \I0/high/ctrlack_internal , 
        \I0/high/nlocalcd , \I0/high/U4/U28/U1/clr , \I0/high/U4/U28/U1/set , 
        \I0/high/U1/Z , \I0/high/U1664/y[0] , \I0/high/U1664/y[1] , 
        \I0/high/U1664/x[1] , \I0/high/U1664/x[3] , \I0/high/U1664/x[2] , 
        \I0/high/U1664/x[0] , \I0/high/U1664/U28/Z , \I0/high/U1664/U32/Z , 
        \I0/high/U1664/U29/Z , \I0/high/U1664/U33/Z , \I0/high/U1664/U30/Z , 
        \I0/high/U1664/U31/Z , \I0/high/U1664/U37/Z , \I0/high/U1669/nr , 
        \I0/high/U1669/nd , \I0/high/U1669/n2 , \I1/net20 , \I1/net33 , 
        \I1/net32 , \I1/low/drivel , \I1/low/driveh , \I1/low/localcd , 
        \I1/low/ncd[7] , \I1/low/ncd[6] , \I1/low/ncd[5] , \I1/low/ncd[4] , 
        \I1/low/ncd[3] , \I1/low/ncd[2] , \I1/low/ncd[1] , \I1/low/ncd[0] , 
        \I1/low/ba , \I1/low/latch , \I1/low/acb , \I1/low/ctrlack_internal , 
        \I1/low/nlocalcd , \I1/low/U4/U28/U1/clr , \I1/low/U4/U28/U1/set , 
        \I1/low/U1/Z , \I1/low/U1664/y[0] , \I1/low/U1664/y[1] , 
        \I1/low/U1664/x[1] , \I1/low/U1664/x[3] , \I1/low/U1664/x[2] , 
        \I1/low/U1664/x[0] , \I1/low/U1664/U28/Z , \I1/low/U1664/U32/Z , 
        \I1/low/U1664/U29/Z , \I1/low/U1664/U33/Z , \I1/low/U1664/U30/Z , 
        \I1/low/U1664/U31/Z , \I1/low/U1664/U37/Z , \I1/low/U1669/nr , 
        \I1/low/U1669/nd , \I1/low/U1669/n2 , \I1/high/drivel , 
        \I1/high/driveh , \I1/high/localcd , \I1/high/ncd[7] , 
        \I1/high/ncd[6] , \I1/high/ncd[5] , \I1/high/ncd[4] , \I1/high/ncd[3] , 
        \I1/high/ncd[2] , \I1/high/ncd[1] , \I1/high/ncd[0] , \I1/high/ba , 
        \I1/high/latch , \I1/high/acb , \I1/high/ctrlack_internal , 
        \I1/high/nlocalcd , \I1/high/U4/U28/U1/clr , \I1/high/U4/U28/U1/set , 
        \I1/high/U1/Z , \I1/high/U1664/y[0] , \I1/high/U1664/y[1] , 
        \I1/high/U1664/x[1] , \I1/high/U1664/x[3] , \I1/high/U1664/x[2] , 
        \I1/high/U1664/x[0] , \I1/high/U1664/U28/Z , \I1/high/U1664/U32/Z , 
        \I1/high/U1664/U29/Z , \I1/high/U1664/U33/Z , \I1/high/U1664/U30/Z , 
        \I1/high/U1664/U31/Z , \I1/high/U1664/U37/Z , \I1/high/U1669/nr , 
        \I1/high/U1669/nd , \I1/high/U1669/n2 , n1, n2, n3, n4, n5, n6, n7, n8;
    nand2_1 \U3/U5  ( .x(pullreq), .a(net30), .b(net31) );
    nor2_1 \I0/U3/U5  ( .x(net30), .a(\I0/net32 ), .b(\I0/net33 ) );
    buf_2 \I0/low/U1653  ( .x(\I0/low/latch ), .a(\I0/net32 ) );
    nor2_1 \I0/low/U264/U5  ( .x(\I0/low/nlocalcd ), .a(reset), .b(
        \I0/low/localcd ) );
    nor2_1 \I0/low/U1659_0_/U5  ( .x(\I0/low/ncd[0] ), .a(ol[0]), .b(oh[0]) );
    nor2_1 \I0/low/U1659_1_/U5  ( .x(\I0/low/ncd[1] ), .a(ol[1]), .b(oh[1]) );
    nor2_1 \I0/low/U1659_2_/U5  ( .x(\I0/low/ncd[2] ), .a(ol[2]), .b(oh[2]) );
    nor2_1 \I0/low/U1659_3_/U5  ( .x(\I0/low/ncd[3] ), .a(ol[3]), .b(oh[3]) );
    nor2_1 \I0/low/U1659_4_/U5  ( .x(\I0/low/ncd[4] ), .a(ol[4]), .b(oh[4]) );
    nor2_1 \I0/low/U1659_5_/U5  ( .x(\I0/low/ncd[5] ), .a(ol[5]), .b(oh[5]) );
    nor2_1 \I0/low/U1659_6_/U5  ( .x(\I0/low/ncd[6] ), .a(ol[6]), .b(oh[6]) );
    nor2_1 \I0/low/U1659_7_/U5  ( .x(\I0/low/ncd[7] ), .a(ol[7]), .b(oh[7]) );
    nor2_1 \I0/low/U3/U5  ( .x(\I0/low/ctrlack_internal ), .a(\I0/low/acb ), 
        .b(\I0/low/ba ) );
    buf_2 \I0/low/U1665/U7  ( .x(\I0/low/driveh ), .a(\I0/net20 ) );
    buf_2 \I0/low/U1666/U7  ( .x(\I0/low/drivel ), .a(\I0/net20 ) );
    ao23_1 \I0/low/U1658_0_/U21/U1/U1  ( .x(ol[0]), .a(\I0/low/driveh ), .b(ol
        [0]), .c(n1), .d(pull_l[0]), .e(n2) );
    ao23_1 \I0/low/U1658_1_/U21/U1/U1  ( .x(ol[1]), .a(\I0/low/drivel ), .b(ol
        [1]), .c(\I0/low/driveh ), .d(pull_l[1]), .e(n2) );
    ao23_1 \I0/low/U1658_2_/U21/U1/U1  ( .x(ol[2]), .a(\I0/low/drivel ), .b(ol
        [2]), .c(\I0/low/driveh ), .d(pull_l[2]), .e(n2) );
    ao23_1 \I0/low/U1658_3_/U21/U1/U1  ( .x(ol[3]), .a(\I0/low/driveh ), .b(ol
        [3]), .c(\I0/low/drivel ), .d(pull_l[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_4_/U21/U1/U1  ( .x(ol[4]), .a(n1), .b(ol[4]), .c(
        \I0/low/drivel ), .d(pull_l[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_5_/U21/U1/U1  ( .x(ol[5]), .a(\I0/low/driveh ), .b(ol
        [5]), .c(n1), .d(pull_l[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_6_/U21/U1/U1  ( .x(ol[6]), .a(\I0/low/drivel ), .b(ol
        [6]), .c(\I0/low/driveh ), .d(pull_l[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_7_/U21/U1/U1  ( .x(ol[7]), .a(n1), .b(ol[7]), .c(n1), 
        .d(pull_l[7]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_0_/U21/U1/U1  ( .x(oh[0]), .a(\I0/low/driveh ), .b(oh
        [0]), .c(n1), .d(pull_h[0]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_1_/U21/U1/U1  ( .x(oh[1]), .a(n1), .b(oh[1]), .c(
        \I0/low/drivel ), .d(pull_h[1]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_2_/U21/U1/U1  ( .x(oh[2]), .a(\I0/low/drivel ), .b(oh
        [2]), .c(\I0/low/drivel ), .d(pull_h[2]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_3_/U21/U1/U1  ( .x(oh[3]), .a(n1), .b(oh[3]), .c(
        \I0/low/driveh ), .d(pull_h[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_4_/U21/U1/U1  ( .x(oh[4]), .a(n1), .b(oh[4]), .c(n1), 
        .d(pull_h[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_5_/U21/U1/U1  ( .x(oh[5]), .a(\I0/low/drivel ), .b(oh
        [5]), .c(n1), .d(pull_h[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_6_/U21/U1/U1  ( .x(oh[6]), .a(\I0/low/drivel ), .b(oh
        [6]), .c(\I0/low/driveh ), .d(pull_h[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_7_/U21/U1/U1  ( .x(oh[7]), .a(\I0/low/driveh ), .b(oh
        [7]), .c(\I0/low/drivel ), .d(pull_h[7]), .e(\I0/low/latch ) );
    aoai211_1 \I0/low/U4/U28/U1/U1  ( .x(\I0/low/U4/U28/U1/clr ), .a(
        \I0/net20 ), .b(\I0/low/acb ), .c(\I0/low/nlocalcd ), .d(\I0/net32 )
         );
    nand3_1 \I0/low/U4/U28/U1/U2  ( .x(\I0/low/U4/U28/U1/set ), .a(
        \I0/low/nlocalcd ), .b(\I0/net20 ), .c(\I0/low/acb ) );
    nand2_2 \I0/low/U4/U28/U1/U3  ( .x(\I0/net32 ), .a(\I0/low/U4/U28/U1/clr ), 
        .b(\I0/low/U4/U28/U1/set ) );
    oai21_1 \I0/low/U1/U30/U1/U1  ( .x(\I0/low/acb ), .a(\I0/low/U1/Z ), .b(
        \I0/low/ba ), .c(\I0/net20 ) );
    inv_1 \I0/low/U1/U30/U1/U2  ( .x(\I0/low/U1/Z ), .a(\I0/low/acb ) );
    ao222_1 \I0/low/U5/U18/U1/U1  ( .x(\I0/low/ba ), .a(\I0/low/latch ), .b(
        pullcd), .c(\I0/low/latch ), .d(\I0/low/ba ), .e(pullcd), .f(
        \I0/low/ba ) );
    aoi222_1 \I0/low/U1664/U28/U30/U1  ( .x(\I0/low/U1664/x[3] ), .a(
        \I0/low/ncd[7] ), .b(\I0/low/ncd[6] ), .c(\I0/low/ncd[7] ), .d(
        \I0/low/U1664/U28/Z ), .e(\I0/low/ncd[6] ), .f(\I0/low/U1664/U28/Z )
         );
    inv_1 \I0/low/U1664/U28/U30/Uinv  ( .x(\I0/low/U1664/U28/Z ), .a(
        \I0/low/U1664/x[3] ) );
    aoi222_1 \I0/low/U1664/U32/U30/U1  ( .x(\I0/low/U1664/x[0] ), .a(
        \I0/low/ncd[1] ), .b(\I0/low/ncd[0] ), .c(\I0/low/ncd[1] ), .d(
        \I0/low/U1664/U32/Z ), .e(\I0/low/ncd[0] ), .f(\I0/low/U1664/U32/Z )
         );
    inv_1 \I0/low/U1664/U32/U30/Uinv  ( .x(\I0/low/U1664/U32/Z ), .a(
        \I0/low/U1664/x[0] ) );
    aoi222_1 \I0/low/U1664/U29/U30/U1  ( .x(\I0/low/U1664/x[2] ), .a(
        \I0/low/ncd[5] ), .b(\I0/low/ncd[4] ), .c(\I0/low/ncd[5] ), .d(
        \I0/low/U1664/U29/Z ), .e(\I0/low/ncd[4] ), .f(\I0/low/U1664/U29/Z )
         );
    inv_1 \I0/low/U1664/U29/U30/Uinv  ( .x(\I0/low/U1664/U29/Z ), .a(
        \I0/low/U1664/x[2] ) );
    aoi222_1 \I0/low/U1664/U33/U30/U1  ( .x(\I0/low/U1664/y[0] ), .a(
        \I0/low/U1664/x[1] ), .b(\I0/low/U1664/x[0] ), .c(\I0/low/U1664/x[1] ), 
        .d(\I0/low/U1664/U33/Z ), .e(\I0/low/U1664/x[0] ), .f(
        \I0/low/U1664/U33/Z ) );
    inv_1 \I0/low/U1664/U33/U30/Uinv  ( .x(\I0/low/U1664/U33/Z ), .a(
        \I0/low/U1664/y[0] ) );
    aoi222_1 \I0/low/U1664/U30/U30/U1  ( .x(\I0/low/U1664/y[1] ), .a(
        \I0/low/U1664/x[3] ), .b(\I0/low/U1664/x[2] ), .c(\I0/low/U1664/x[3] ), 
        .d(\I0/low/U1664/U30/Z ), .e(\I0/low/U1664/x[2] ), .f(
        \I0/low/U1664/U30/Z ) );
    inv_1 \I0/low/U1664/U30/U30/Uinv  ( .x(\I0/low/U1664/U30/Z ), .a(
        \I0/low/U1664/y[1] ) );
    aoi222_1 \I0/low/U1664/U31/U30/U1  ( .x(\I0/low/U1664/x[1] ), .a(
        \I0/low/ncd[3] ), .b(\I0/low/ncd[2] ), .c(\I0/low/ncd[3] ), .d(
        \I0/low/U1664/U31/Z ), .e(\I0/low/ncd[2] ), .f(\I0/low/U1664/U31/Z )
         );
    inv_1 \I0/low/U1664/U31/U30/Uinv  ( .x(\I0/low/U1664/U31/Z ), .a(
        \I0/low/U1664/x[1] ) );
    aoi222_1 \I0/low/U1664/U37/U30/U1  ( .x(\I0/low/localcd ), .a(
        \I0/low/U1664/y[0] ), .b(\I0/low/U1664/y[1] ), .c(\I0/low/U1664/y[0] ), 
        .d(\I0/low/U1664/U37/Z ), .e(\I0/low/U1664/y[1] ), .f(
        \I0/low/U1664/U37/Z ) );
    inv_1 \I0/low/U1664/U37/U30/Uinv  ( .x(\I0/low/U1664/U37/Z ), .a(
        \I0/low/localcd ) );
    nor3_1 \I0/low/U1669/Unr  ( .x(\I0/low/U1669/nr ), .a(
        \I0/low/ctrlack_internal ), .b(n1), .c(\I0/low/driveh ) );
    nand3_1 \I0/low/U1669/Und  ( .x(\I0/low/U1669/nd ), .a(
        \I0/low/ctrlack_internal ), .b(\I0/low/drivel ), .c(\I0/low/driveh )
         );
    oa21_1 \I0/low/U1669/U1  ( .x(\I0/low/U1669/n2 ), .a(\I0/low/U1669/n2 ), 
        .b(\I0/low/U1669/nr ), .c(\I0/low/U1669/nd ) );
    inv_2 \I0/low/U1669/U3  ( .x(ctrlack), .a(\I0/low/U1669/n2 ) );
    buf_2 \I0/high/U1653  ( .x(\I0/high/latch ), .a(\I0/net33 ) );
    nor2_1 \I0/high/U264/U5  ( .x(\I0/high/nlocalcd ), .a(reset), .b(
        \I0/high/localcd ) );
    nor2_1 \I0/high/U1659_0_/U5  ( .x(\I0/high/ncd[0] ), .a(ol[8]), .b(oh[8])
         );
    nor2_1 \I0/high/U1659_1_/U5  ( .x(\I0/high/ncd[1] ), .a(ol[9]), .b(oh[9])
         );
    nor2_1 \I0/high/U1659_2_/U5  ( .x(\I0/high/ncd[2] ), .a(ol[10]), .b(oh[10]
        ) );
    nor2_1 \I0/high/U1659_3_/U5  ( .x(\I0/high/ncd[3] ), .a(ol[11]), .b(oh[11]
        ) );
    nor2_1 \I0/high/U1659_4_/U5  ( .x(\I0/high/ncd[4] ), .a(ol[12]), .b(oh[12]
        ) );
    nor2_1 \I0/high/U1659_5_/U5  ( .x(\I0/high/ncd[5] ), .a(ol[13]), .b(oh[13]
        ) );
    nor2_1 \I0/high/U1659_6_/U5  ( .x(\I0/high/ncd[6] ), .a(ol[14]), .b(oh[14]
        ) );
    nor2_1 \I0/high/U1659_7_/U5  ( .x(\I0/high/ncd[7] ), .a(ol[15]), .b(oh[15]
        ) );
    nor2_1 \I0/high/U3/U5  ( .x(\I0/high/ctrlack_internal ), .a(\I0/high/acb ), 
        .b(\I0/high/ba ) );
    buf_2 \I0/high/U1665/U7  ( .x(\I0/high/driveh ), .a(net17) );
    buf_2 \I0/high/U1666/U7  ( .x(\I0/high/drivel ), .a(net17) );
    ao23_1 \I0/high/U1658_0_/U21/U1/U1  ( .x(ol[8]), .a(\I0/high/driveh ), .b(
        ol[8]), .c(n3), .d(pull_l[0]), .e(n4) );
    ao23_1 \I0/high/U1658_1_/U21/U1/U1  ( .x(ol[9]), .a(\I0/high/drivel ), .b(
        ol[9]), .c(\I0/high/driveh ), .d(pull_l[1]), .e(n4) );
    ao23_1 \I0/high/U1658_2_/U21/U1/U1  ( .x(ol[10]), .a(\I0/high/drivel ), 
        .b(ol[10]), .c(\I0/high/driveh ), .d(pull_l[2]), .e(n4) );
    ao23_1 \I0/high/U1658_3_/U21/U1/U1  ( .x(ol[11]), .a(\I0/high/driveh ), 
        .b(ol[11]), .c(\I0/high/drivel ), .d(pull_l[3]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_4_/U21/U1/U1  ( .x(ol[12]), .a(n3), .b(ol[12]), .c(
        \I0/high/drivel ), .d(pull_l[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_5_/U21/U1/U1  ( .x(ol[13]), .a(\I0/high/driveh ), 
        .b(ol[13]), .c(n3), .d(pull_l[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_6_/U21/U1/U1  ( .x(ol[14]), .a(\I0/high/drivel ), 
        .b(ol[14]), .c(\I0/high/driveh ), .d(pull_l[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_7_/U21/U1/U1  ( .x(ol[15]), .a(n3), .b(ol[15]), .c(
        n3), .d(pull_l[7]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_0_/U21/U1/U1  ( .x(oh[8]), .a(\I0/high/driveh ), .b(
        oh[8]), .c(n3), .d(pull_h[0]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_1_/U21/U1/U1  ( .x(oh[9]), .a(n3), .b(oh[9]), .c(
        \I0/high/drivel ), .d(pull_h[1]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_2_/U21/U1/U1  ( .x(oh[10]), .a(\I0/high/drivel ), 
        .b(oh[10]), .c(\I0/high/drivel ), .d(pull_h[2]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_3_/U21/U1/U1  ( .x(oh[11]), .a(n3), .b(oh[11]), .c(
        \I0/high/driveh ), .d(pull_h[3]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_4_/U21/U1/U1  ( .x(oh[12]), .a(n3), .b(oh[12]), .c(
        n3), .d(pull_h[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_5_/U21/U1/U1  ( .x(oh[13]), .a(\I0/high/drivel ), 
        .b(oh[13]), .c(n3), .d(pull_h[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_6_/U21/U1/U1  ( .x(oh[14]), .a(\I0/high/drivel ), 
        .b(oh[14]), .c(\I0/high/driveh ), .d(pull_h[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_7_/U21/U1/U1  ( .x(oh[15]), .a(\I0/high/driveh ), 
        .b(oh[15]), .c(\I0/high/drivel ), .d(pull_h[7]), .e(\I0/high/latch )
         );
    aoai211_1 \I0/high/U4/U28/U1/U1  ( .x(\I0/high/U4/U28/U1/clr ), .a(net17), 
        .b(\I0/high/acb ), .c(\I0/high/nlocalcd ), .d(\I0/net33 ) );
    nand3_1 \I0/high/U4/U28/U1/U2  ( .x(\I0/high/U4/U28/U1/set ), .a(
        \I0/high/nlocalcd ), .b(net17), .c(\I0/high/acb ) );
    nand2_2 \I0/high/U4/U28/U1/U3  ( .x(\I0/net33 ), .a(
        \I0/high/U4/U28/U1/clr ), .b(\I0/high/U4/U28/U1/set ) );
    oai21_1 \I0/high/U1/U30/U1/U1  ( .x(\I0/high/acb ), .a(\I0/high/U1/Z ), 
        .b(\I0/high/ba ), .c(net17) );
    inv_1 \I0/high/U1/U30/U1/U2  ( .x(\I0/high/U1/Z ), .a(\I0/high/acb ) );
    ao222_1 \I0/high/U5/U18/U1/U1  ( .x(\I0/high/ba ), .a(\I0/high/latch ), 
        .b(pullcd), .c(\I0/high/latch ), .d(\I0/high/ba ), .e(pullcd), .f(
        \I0/high/ba ) );
    aoi222_1 \I0/high/U1664/U28/U30/U1  ( .x(\I0/high/U1664/x[3] ), .a(
        \I0/high/ncd[7] ), .b(\I0/high/ncd[6] ), .c(\I0/high/ncd[7] ), .d(
        \I0/high/U1664/U28/Z ), .e(\I0/high/ncd[6] ), .f(\I0/high/U1664/U28/Z 
        ) );
    inv_1 \I0/high/U1664/U28/U30/Uinv  ( .x(\I0/high/U1664/U28/Z ), .a(
        \I0/high/U1664/x[3] ) );
    aoi222_1 \I0/high/U1664/U32/U30/U1  ( .x(\I0/high/U1664/x[0] ), .a(
        \I0/high/ncd[1] ), .b(\I0/high/ncd[0] ), .c(\I0/high/ncd[1] ), .d(
        \I0/high/U1664/U32/Z ), .e(\I0/high/ncd[0] ), .f(\I0/high/U1664/U32/Z 
        ) );
    inv_1 \I0/high/U1664/U32/U30/Uinv  ( .x(\I0/high/U1664/U32/Z ), .a(
        \I0/high/U1664/x[0] ) );
    aoi222_1 \I0/high/U1664/U29/U30/U1  ( .x(\I0/high/U1664/x[2] ), .a(
        \I0/high/ncd[5] ), .b(\I0/high/ncd[4] ), .c(\I0/high/ncd[5] ), .d(
        \I0/high/U1664/U29/Z ), .e(\I0/high/ncd[4] ), .f(\I0/high/U1664/U29/Z 
        ) );
    inv_1 \I0/high/U1664/U29/U30/Uinv  ( .x(\I0/high/U1664/U29/Z ), .a(
        \I0/high/U1664/x[2] ) );
    aoi222_1 \I0/high/U1664/U33/U30/U1  ( .x(\I0/high/U1664/y[0] ), .a(
        \I0/high/U1664/x[1] ), .b(\I0/high/U1664/x[0] ), .c(
        \I0/high/U1664/x[1] ), .d(\I0/high/U1664/U33/Z ), .e(
        \I0/high/U1664/x[0] ), .f(\I0/high/U1664/U33/Z ) );
    inv_1 \I0/high/U1664/U33/U30/Uinv  ( .x(\I0/high/U1664/U33/Z ), .a(
        \I0/high/U1664/y[0] ) );
    aoi222_1 \I0/high/U1664/U30/U30/U1  ( .x(\I0/high/U1664/y[1] ), .a(
        \I0/high/U1664/x[3] ), .b(\I0/high/U1664/x[2] ), .c(
        \I0/high/U1664/x[3] ), .d(\I0/high/U1664/U30/Z ), .e(
        \I0/high/U1664/x[2] ), .f(\I0/high/U1664/U30/Z ) );
    inv_1 \I0/high/U1664/U30/U30/Uinv  ( .x(\I0/high/U1664/U30/Z ), .a(
        \I0/high/U1664/y[1] ) );
    aoi222_1 \I0/high/U1664/U31/U30/U1  ( .x(\I0/high/U1664/x[1] ), .a(
        \I0/high/ncd[3] ), .b(\I0/high/ncd[2] ), .c(\I0/high/ncd[3] ), .d(
        \I0/high/U1664/U31/Z ), .e(\I0/high/ncd[2] ), .f(\I0/high/U1664/U31/Z 
        ) );
    inv_1 \I0/high/U1664/U31/U30/Uinv  ( .x(\I0/high/U1664/U31/Z ), .a(
        \I0/high/U1664/x[1] ) );
    aoi222_1 \I0/high/U1664/U37/U30/U1  ( .x(\I0/high/localcd ), .a(
        \I0/high/U1664/y[0] ), .b(\I0/high/U1664/y[1] ), .c(
        \I0/high/U1664/y[0] ), .d(\I0/high/U1664/U37/Z ), .e(
        \I0/high/U1664/y[1] ), .f(\I0/high/U1664/U37/Z ) );
    inv_1 \I0/high/U1664/U37/U30/Uinv  ( .x(\I0/high/U1664/U37/Z ), .a(
        \I0/high/localcd ) );
    nor3_1 \I0/high/U1669/Unr  ( .x(\I0/high/U1669/nr ), .a(
        \I0/high/ctrlack_internal ), .b(n3), .c(\I0/high/driveh ) );
    nand3_1 \I0/high/U1669/Und  ( .x(\I0/high/U1669/nd ), .a(
        \I0/high/ctrlack_internal ), .b(\I0/high/drivel ), .c(\I0/high/driveh 
        ) );
    oa21_1 \I0/high/U1669/U1  ( .x(\I0/high/U1669/n2 ), .a(\I0/high/U1669/n2 ), 
        .b(\I0/high/U1669/nr ), .c(\I0/high/U1669/nd ) );
    inv_2 \I0/high/U1669/U3  ( .x(\I0/net20 ), .a(\I0/high/U1669/n2 ) );
    nor2_1 \I1/U3/U5  ( .x(net31), .a(\I1/net32 ), .b(\I1/net33 ) );
    buf_2 \I1/low/U1653  ( .x(\I1/low/latch ), .a(\I1/net32 ) );
    nor2_1 \I1/low/U264/U5  ( .x(\I1/low/nlocalcd ), .a(reset), .b(
        \I1/low/localcd ) );
    nor2_1 \I1/low/U1659_0_/U5  ( .x(\I1/low/ncd[0] ), .a(ol[16]), .b(oh[16])
         );
    nor2_1 \I1/low/U1659_1_/U5  ( .x(\I1/low/ncd[1] ), .a(ol[17]), .b(oh[17])
         );
    nor2_1 \I1/low/U1659_2_/U5  ( .x(\I1/low/ncd[2] ), .a(ol[18]), .b(oh[18])
         );
    nor2_1 \I1/low/U1659_3_/U5  ( .x(\I1/low/ncd[3] ), .a(ol[19]), .b(oh[19])
         );
    nor2_1 \I1/low/U1659_4_/U5  ( .x(\I1/low/ncd[4] ), .a(ol[20]), .b(oh[20])
         );
    nor2_1 \I1/low/U1659_5_/U5  ( .x(\I1/low/ncd[5] ), .a(ol[21]), .b(oh[21])
         );
    nor2_1 \I1/low/U1659_6_/U5  ( .x(\I1/low/ncd[6] ), .a(ol[22]), .b(oh[22])
         );
    nor2_1 \I1/low/U1659_7_/U5  ( .x(\I1/low/ncd[7] ), .a(ol[23]), .b(oh[23])
         );
    nor2_1 \I1/low/U3/U5  ( .x(\I1/low/ctrlack_internal ), .a(\I1/low/acb ), 
        .b(\I1/low/ba ) );
    buf_2 \I1/low/U1665/U7  ( .x(\I1/low/driveh ), .a(\I1/net20 ) );
    buf_2 \I1/low/U1666/U7  ( .x(\I1/low/drivel ), .a(\I1/net20 ) );
    ao23_1 \I1/low/U1658_0_/U21/U1/U1  ( .x(ol[16]), .a(\I1/low/driveh ), .b(
        ol[16]), .c(n5), .d(pull_l[0]), .e(n6) );
    ao23_1 \I1/low/U1658_1_/U21/U1/U1  ( .x(ol[17]), .a(\I1/low/drivel ), .b(
        ol[17]), .c(\I1/low/driveh ), .d(pull_l[1]), .e(n6) );
    ao23_1 \I1/low/U1658_2_/U21/U1/U1  ( .x(ol[18]), .a(\I1/low/drivel ), .b(
        ol[18]), .c(\I1/low/driveh ), .d(pull_l[2]), .e(n6) );
    ao23_1 \I1/low/U1658_3_/U21/U1/U1  ( .x(ol[19]), .a(\I1/low/driveh ), .b(
        ol[19]), .c(\I1/low/drivel ), .d(pull_l[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_4_/U21/U1/U1  ( .x(ol[20]), .a(n5), .b(ol[20]), .c(
        \I1/low/drivel ), .d(pull_l[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_5_/U21/U1/U1  ( .x(ol[21]), .a(\I1/low/driveh ), .b(
        ol[21]), .c(n5), .d(pull_l[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_6_/U21/U1/U1  ( .x(ol[22]), .a(\I1/low/drivel ), .b(
        ol[22]), .c(\I1/low/driveh ), .d(pull_l[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_7_/U21/U1/U1  ( .x(ol[23]), .a(n5), .b(ol[23]), .c(n5
        ), .d(pull_l[7]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_0_/U21/U1/U1  ( .x(oh[16]), .a(\I1/low/driveh ), .b(
        oh[16]), .c(n5), .d(pull_h[0]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_1_/U21/U1/U1  ( .x(oh[17]), .a(n5), .b(oh[17]), .c(
        \I1/low/drivel ), .d(pull_h[1]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_2_/U21/U1/U1  ( .x(oh[18]), .a(\I1/low/drivel ), .b(
        oh[18]), .c(\I1/low/drivel ), .d(pull_h[2]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_3_/U21/U1/U1  ( .x(oh[19]), .a(n5), .b(oh[19]), .c(
        \I1/low/driveh ), .d(pull_h[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_4_/U21/U1/U1  ( .x(oh[20]), .a(n5), .b(oh[20]), .c(n5
        ), .d(pull_h[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_5_/U21/U1/U1  ( .x(oh[21]), .a(\I1/low/drivel ), .b(
        oh[21]), .c(n5), .d(pull_h[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_6_/U21/U1/U1  ( .x(oh[22]), .a(\I1/low/drivel ), .b(
        oh[22]), .c(\I1/low/driveh ), .d(pull_h[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_7_/U21/U1/U1  ( .x(oh[23]), .a(\I1/low/driveh ), .b(
        oh[23]), .c(\I1/low/drivel ), .d(pull_h[7]), .e(\I1/low/latch ) );
    aoai211_1 \I1/low/U4/U28/U1/U1  ( .x(\I1/low/U4/U28/U1/clr ), .a(
        \I1/net20 ), .b(\I1/low/acb ), .c(\I1/low/nlocalcd ), .d(\I1/net32 )
         );
    nand3_1 \I1/low/U4/U28/U1/U2  ( .x(\I1/low/U4/U28/U1/set ), .a(
        \I1/low/nlocalcd ), .b(\I1/net20 ), .c(\I1/low/acb ) );
    nand2_2 \I1/low/U4/U28/U1/U3  ( .x(\I1/net32 ), .a(\I1/low/U4/U28/U1/clr ), 
        .b(\I1/low/U4/U28/U1/set ) );
    oai21_1 \I1/low/U1/U30/U1/U1  ( .x(\I1/low/acb ), .a(\I1/low/U1/Z ), .b(
        \I1/low/ba ), .c(\I1/net20 ) );
    inv_1 \I1/low/U1/U30/U1/U2  ( .x(\I1/low/U1/Z ), .a(\I1/low/acb ) );
    ao222_1 \I1/low/U5/U18/U1/U1  ( .x(\I1/low/ba ), .a(\I1/low/latch ), .b(
        pullcd), .c(\I1/low/latch ), .d(\I1/low/ba ), .e(pullcd), .f(
        \I1/low/ba ) );
    aoi222_1 \I1/low/U1664/U28/U30/U1  ( .x(\I1/low/U1664/x[3] ), .a(
        \I1/low/ncd[7] ), .b(\I1/low/ncd[6] ), .c(\I1/low/ncd[7] ), .d(
        \I1/low/U1664/U28/Z ), .e(\I1/low/ncd[6] ), .f(\I1/low/U1664/U28/Z )
         );
    inv_1 \I1/low/U1664/U28/U30/Uinv  ( .x(\I1/low/U1664/U28/Z ), .a(
        \I1/low/U1664/x[3] ) );
    aoi222_1 \I1/low/U1664/U32/U30/U1  ( .x(\I1/low/U1664/x[0] ), .a(
        \I1/low/ncd[1] ), .b(\I1/low/ncd[0] ), .c(\I1/low/ncd[1] ), .d(
        \I1/low/U1664/U32/Z ), .e(\I1/low/ncd[0] ), .f(\I1/low/U1664/U32/Z )
         );
    inv_1 \I1/low/U1664/U32/U30/Uinv  ( .x(\I1/low/U1664/U32/Z ), .a(
        \I1/low/U1664/x[0] ) );
    aoi222_1 \I1/low/U1664/U29/U30/U1  ( .x(\I1/low/U1664/x[2] ), .a(
        \I1/low/ncd[5] ), .b(\I1/low/ncd[4] ), .c(\I1/low/ncd[5] ), .d(
        \I1/low/U1664/U29/Z ), .e(\I1/low/ncd[4] ), .f(\I1/low/U1664/U29/Z )
         );
    inv_1 \I1/low/U1664/U29/U30/Uinv  ( .x(\I1/low/U1664/U29/Z ), .a(
        \I1/low/U1664/x[2] ) );
    aoi222_1 \I1/low/U1664/U33/U30/U1  ( .x(\I1/low/U1664/y[0] ), .a(
        \I1/low/U1664/x[1] ), .b(\I1/low/U1664/x[0] ), .c(\I1/low/U1664/x[1] ), 
        .d(\I1/low/U1664/U33/Z ), .e(\I1/low/U1664/x[0] ), .f(
        \I1/low/U1664/U33/Z ) );
    inv_1 \I1/low/U1664/U33/U30/Uinv  ( .x(\I1/low/U1664/U33/Z ), .a(
        \I1/low/U1664/y[0] ) );
    aoi222_1 \I1/low/U1664/U30/U30/U1  ( .x(\I1/low/U1664/y[1] ), .a(
        \I1/low/U1664/x[3] ), .b(\I1/low/U1664/x[2] ), .c(\I1/low/U1664/x[3] ), 
        .d(\I1/low/U1664/U30/Z ), .e(\I1/low/U1664/x[2] ), .f(
        \I1/low/U1664/U30/Z ) );
    inv_1 \I1/low/U1664/U30/U30/Uinv  ( .x(\I1/low/U1664/U30/Z ), .a(
        \I1/low/U1664/y[1] ) );
    aoi222_1 \I1/low/U1664/U31/U30/U1  ( .x(\I1/low/U1664/x[1] ), .a(
        \I1/low/ncd[3] ), .b(\I1/low/ncd[2] ), .c(\I1/low/ncd[3] ), .d(
        \I1/low/U1664/U31/Z ), .e(\I1/low/ncd[2] ), .f(\I1/low/U1664/U31/Z )
         );
    inv_1 \I1/low/U1664/U31/U30/Uinv  ( .x(\I1/low/U1664/U31/Z ), .a(
        \I1/low/U1664/x[1] ) );
    aoi222_1 \I1/low/U1664/U37/U30/U1  ( .x(\I1/low/localcd ), .a(
        \I1/low/U1664/y[0] ), .b(\I1/low/U1664/y[1] ), .c(\I1/low/U1664/y[0] ), 
        .d(\I1/low/U1664/U37/Z ), .e(\I1/low/U1664/y[1] ), .f(
        \I1/low/U1664/U37/Z ) );
    inv_1 \I1/low/U1664/U37/U30/Uinv  ( .x(\I1/low/U1664/U37/Z ), .a(
        \I1/low/localcd ) );
    nor3_1 \I1/low/U1669/Unr  ( .x(\I1/low/U1669/nr ), .a(
        \I1/low/ctrlack_internal ), .b(n5), .c(\I1/low/driveh ) );
    nand3_1 \I1/low/U1669/Und  ( .x(\I1/low/U1669/nd ), .a(
        \I1/low/ctrlack_internal ), .b(\I1/low/drivel ), .c(\I1/low/driveh )
         );
    oa21_1 \I1/low/U1669/U1  ( .x(\I1/low/U1669/n2 ), .a(\I1/low/U1669/n2 ), 
        .b(\I1/low/U1669/nr ), .c(\I1/low/U1669/nd ) );
    inv_2 \I1/low/U1669/U3  ( .x(net17), .a(\I1/low/U1669/n2 ) );
    buf_2 \I1/high/U1653  ( .x(\I1/high/latch ), .a(\I1/net33 ) );
    nor2_1 \I1/high/U264/U5  ( .x(\I1/high/nlocalcd ), .a(reset), .b(
        \I1/high/localcd ) );
    nor2_1 \I1/high/U1659_0_/U5  ( .x(\I1/high/ncd[0] ), .a(ol[24]), .b(oh[24]
        ) );
    nor2_1 \I1/high/U1659_1_/U5  ( .x(\I1/high/ncd[1] ), .a(ol[25]), .b(oh[25]
        ) );
    nor2_1 \I1/high/U1659_2_/U5  ( .x(\I1/high/ncd[2] ), .a(ol[26]), .b(oh[26]
        ) );
    nor2_1 \I1/high/U1659_3_/U5  ( .x(\I1/high/ncd[3] ), .a(ol[27]), .b(oh[27]
        ) );
    nor2_1 \I1/high/U1659_4_/U5  ( .x(\I1/high/ncd[4] ), .a(ol[28]), .b(oh[28]
        ) );
    nor2_1 \I1/high/U1659_5_/U5  ( .x(\I1/high/ncd[5] ), .a(ol[29]), .b(oh[29]
        ) );
    nor2_1 \I1/high/U1659_6_/U5  ( .x(\I1/high/ncd[6] ), .a(ol[30]), .b(oh[30]
        ) );
    nor2_1 \I1/high/U1659_7_/U5  ( .x(\I1/high/ncd[7] ), .a(ol[31]), .b(oh[31]
        ) );
    nor2_1 \I1/high/U3/U5  ( .x(\I1/high/ctrlack_internal ), .a(\I1/high/acb ), 
        .b(\I1/high/ba ) );
    buf_2 \I1/high/U1665/U7  ( .x(\I1/high/driveh ), .a(ctrlreq) );
    buf_2 \I1/high/U1666/U7  ( .x(\I1/high/drivel ), .a(ctrlreq) );
    ao23_1 \I1/high/U1658_0_/U21/U1/U1  ( .x(ol[24]), .a(\I1/high/driveh ), 
        .b(ol[24]), .c(n7), .d(pull_l[0]), .e(n8) );
    ao23_1 \I1/high/U1658_1_/U21/U1/U1  ( .x(ol[25]), .a(\I1/high/drivel ), 
        .b(ol[25]), .c(\I1/high/driveh ), .d(pull_l[1]), .e(n8) );
    ao23_1 \I1/high/U1658_2_/U21/U1/U1  ( .x(ol[26]), .a(\I1/high/drivel ), 
        .b(ol[26]), .c(\I1/high/driveh ), .d(pull_l[2]), .e(n8) );
    ao23_1 \I1/high/U1658_3_/U21/U1/U1  ( .x(ol[27]), .a(\I1/high/driveh ), 
        .b(ol[27]), .c(\I1/high/drivel ), .d(pull_l[3]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1658_4_/U21/U1/U1  ( .x(ol[28]), .a(n7), .b(ol[28]), .c(
        \I1/high/drivel ), .d(pull_l[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_5_/U21/U1/U1  ( .x(ol[29]), .a(\I1/high/driveh ), 
        .b(ol[29]), .c(n7), .d(pull_l[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_6_/U21/U1/U1  ( .x(ol[30]), .a(\I1/high/drivel ), 
        .b(ol[30]), .c(\I1/high/driveh ), .d(pull_l[6]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1658_7_/U21/U1/U1  ( .x(ol[31]), .a(n7), .b(ol[31]), .c(
        n7), .d(pull_l[7]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_0_/U21/U1/U1  ( .x(oh[24]), .a(\I1/high/driveh ), 
        .b(oh[24]), .c(n7), .d(pull_h[0]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_1_/U21/U1/U1  ( .x(oh[25]), .a(n7), .b(oh[25]), .c(
        \I1/high/drivel ), .d(pull_h[1]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_2_/U21/U1/U1  ( .x(oh[26]), .a(\I1/high/drivel ), 
        .b(oh[26]), .c(\I1/high/drivel ), .d(pull_h[2]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1651_3_/U21/U1/U1  ( .x(oh[27]), .a(n7), .b(oh[27]), .c(
        \I1/high/driveh ), .d(pull_h[3]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_4_/U21/U1/U1  ( .x(oh[28]), .a(n7), .b(oh[28]), .c(
        n7), .d(pull_h[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_5_/U21/U1/U1  ( .x(oh[29]), .a(\I1/high/drivel ), 
        .b(oh[29]), .c(n7), .d(pull_h[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_6_/U21/U1/U1  ( .x(oh[30]), .a(\I1/high/drivel ), 
        .b(oh[30]), .c(\I1/high/driveh ), .d(pull_h[6]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1651_7_/U21/U1/U1  ( .x(oh[31]), .a(\I1/high/driveh ), 
        .b(oh[31]), .c(\I1/high/drivel ), .d(pull_h[7]), .e(\I1/high/latch )
         );
    aoai211_1 \I1/high/U4/U28/U1/U1  ( .x(\I1/high/U4/U28/U1/clr ), .a(ctrlreq
        ), .b(\I1/high/acb ), .c(\I1/high/nlocalcd ), .d(\I1/net33 ) );
    nand3_1 \I1/high/U4/U28/U1/U2  ( .x(\I1/high/U4/U28/U1/set ), .a(
        \I1/high/nlocalcd ), .b(ctrlreq), .c(\I1/high/acb ) );
    nand2_2 \I1/high/U4/U28/U1/U3  ( .x(\I1/net33 ), .a(
        \I1/high/U4/U28/U1/clr ), .b(\I1/high/U4/U28/U1/set ) );
    oai21_1 \I1/high/U1/U30/U1/U1  ( .x(\I1/high/acb ), .a(\I1/high/U1/Z ), 
        .b(\I1/high/ba ), .c(ctrlreq) );
    inv_1 \I1/high/U1/U30/U1/U2  ( .x(\I1/high/U1/Z ), .a(\I1/high/acb ) );
    ao222_1 \I1/high/U5/U18/U1/U1  ( .x(\I1/high/ba ), .a(\I1/high/latch ), 
        .b(pullcd), .c(\I1/high/latch ), .d(\I1/high/ba ), .e(pullcd), .f(
        \I1/high/ba ) );
    aoi222_1 \I1/high/U1664/U28/U30/U1  ( .x(\I1/high/U1664/x[3] ), .a(
        \I1/high/ncd[7] ), .b(\I1/high/ncd[6] ), .c(\I1/high/ncd[7] ), .d(
        \I1/high/U1664/U28/Z ), .e(\I1/high/ncd[6] ), .f(\I1/high/U1664/U28/Z 
        ) );
    inv_1 \I1/high/U1664/U28/U30/Uinv  ( .x(\I1/high/U1664/U28/Z ), .a(
        \I1/high/U1664/x[3] ) );
    aoi222_1 \I1/high/U1664/U32/U30/U1  ( .x(\I1/high/U1664/x[0] ), .a(
        \I1/high/ncd[1] ), .b(\I1/high/ncd[0] ), .c(\I1/high/ncd[1] ), .d(
        \I1/high/U1664/U32/Z ), .e(\I1/high/ncd[0] ), .f(\I1/high/U1664/U32/Z 
        ) );
    inv_1 \I1/high/U1664/U32/U30/Uinv  ( .x(\I1/high/U1664/U32/Z ), .a(
        \I1/high/U1664/x[0] ) );
    aoi222_1 \I1/high/U1664/U29/U30/U1  ( .x(\I1/high/U1664/x[2] ), .a(
        \I1/high/ncd[5] ), .b(\I1/high/ncd[4] ), .c(\I1/high/ncd[5] ), .d(
        \I1/high/U1664/U29/Z ), .e(\I1/high/ncd[4] ), .f(\I1/high/U1664/U29/Z 
        ) );
    inv_1 \I1/high/U1664/U29/U30/Uinv  ( .x(\I1/high/U1664/U29/Z ), .a(
        \I1/high/U1664/x[2] ) );
    aoi222_1 \I1/high/U1664/U33/U30/U1  ( .x(\I1/high/U1664/y[0] ), .a(
        \I1/high/U1664/x[1] ), .b(\I1/high/U1664/x[0] ), .c(
        \I1/high/U1664/x[1] ), .d(\I1/high/U1664/U33/Z ), .e(
        \I1/high/U1664/x[0] ), .f(\I1/high/U1664/U33/Z ) );
    inv_1 \I1/high/U1664/U33/U30/Uinv  ( .x(\I1/high/U1664/U33/Z ), .a(
        \I1/high/U1664/y[0] ) );
    aoi222_1 \I1/high/U1664/U30/U30/U1  ( .x(\I1/high/U1664/y[1] ), .a(
        \I1/high/U1664/x[3] ), .b(\I1/high/U1664/x[2] ), .c(
        \I1/high/U1664/x[3] ), .d(\I1/high/U1664/U30/Z ), .e(
        \I1/high/U1664/x[2] ), .f(\I1/high/U1664/U30/Z ) );
    inv_1 \I1/high/U1664/U30/U30/Uinv  ( .x(\I1/high/U1664/U30/Z ), .a(
        \I1/high/U1664/y[1] ) );
    aoi222_1 \I1/high/U1664/U31/U30/U1  ( .x(\I1/high/U1664/x[1] ), .a(
        \I1/high/ncd[3] ), .b(\I1/high/ncd[2] ), .c(\I1/high/ncd[3] ), .d(
        \I1/high/U1664/U31/Z ), .e(\I1/high/ncd[2] ), .f(\I1/high/U1664/U31/Z 
        ) );
    inv_1 \I1/high/U1664/U31/U30/Uinv  ( .x(\I1/high/U1664/U31/Z ), .a(
        \I1/high/U1664/x[1] ) );
    aoi222_1 \I1/high/U1664/U37/U30/U1  ( .x(\I1/high/localcd ), .a(
        \I1/high/U1664/y[0] ), .b(\I1/high/U1664/y[1] ), .c(
        \I1/high/U1664/y[0] ), .d(\I1/high/U1664/U37/Z ), .e(
        \I1/high/U1664/y[1] ), .f(\I1/high/U1664/U37/Z ) );
    inv_1 \I1/high/U1664/U37/U30/Uinv  ( .x(\I1/high/U1664/U37/Z ), .a(
        \I1/high/localcd ) );
    nor3_1 \I1/high/U1669/Unr  ( .x(\I1/high/U1669/nr ), .a(
        \I1/high/ctrlack_internal ), .b(n7), .c(\I1/high/driveh ) );
    nand3_1 \I1/high/U1669/Und  ( .x(\I1/high/U1669/nd ), .a(
        \I1/high/ctrlack_internal ), .b(\I1/high/drivel ), .c(\I1/high/driveh 
        ) );
    oa21_1 \I1/high/U1669/U1  ( .x(\I1/high/U1669/n2 ), .a(\I1/high/U1669/n2 ), 
        .b(\I1/high/U1669/nr ), .c(\I1/high/U1669/nd ) );
    inv_2 \I1/high/U1669/U3  ( .x(\I1/net20 ), .a(\I1/high/U1669/n2 ) );
    buf_2 U1 ( .x(n1), .a(\I0/net20 ) );
    buf_1 U2 ( .x(n2), .a(\I0/low/latch ) );
    buf_2 U3 ( .x(n3), .a(net17) );
    buf_1 U4 ( .x(n4), .a(\I0/high/latch ) );
    buf_2 U5 ( .x(n5), .a(\I1/net20 ) );
    buf_1 U6 ( .x(n6), .a(\I1/low/latch ) );
    buf_2 U7 ( .x(n7), .a(ctrlreq) );
    buf_1 U8 ( .x(n8), .a(\I1/high/latch ) );
endmodule


module chain_irdemux_32new_5 ( ctrlack, oh, ol, pullreq, pull_h, pull_l, 
    pullcd, reset, ctrlreq );
output [31:0] oh;
output [31:0] ol;
input  [7:0] pull_h;
input  [7:0] pull_l;
input  pullcd, reset, ctrlreq;
output ctrlack, pullreq;
    wire net30, net31, net17, \I0/net20 , \I0/net33 , \I0/net32 , 
        \I0/low/drivel , \I0/low/driveh , \I0/low/localcd , \I0/low/ncd[7] , 
        \I0/low/ncd[6] , \I0/low/ncd[5] , \I0/low/ncd[4] , \I0/low/ncd[3] , 
        \I0/low/ncd[2] , \I0/low/ncd[1] , \I0/low/ncd[0] , \I0/low/ba , 
        \I0/low/latch , \I0/low/acb , \I0/low/ctrlack_internal , 
        \I0/low/nlocalcd , \I0/low/U4/U28/U1/clr , \I0/low/U4/U28/U1/set , 
        \I0/low/U1/Z , \I0/low/U1664/y[0] , \I0/low/U1664/y[1] , 
        \I0/low/U1664/x[1] , \I0/low/U1664/x[3] , \I0/low/U1664/x[2] , 
        \I0/low/U1664/x[0] , \I0/low/U1664/U28/Z , \I0/low/U1664/U32/Z , 
        \I0/low/U1664/U29/Z , \I0/low/U1664/U33/Z , \I0/low/U1664/U30/Z , 
        \I0/low/U1664/U31/Z , \I0/low/U1664/U37/Z , \I0/low/U1669/nr , 
        \I0/low/U1669/nd , \I0/low/U1669/n2 , \I0/high/drivel , 
        \I0/high/driveh , \I0/high/localcd , \I0/high/ncd[7] , 
        \I0/high/ncd[6] , \I0/high/ncd[5] , \I0/high/ncd[4] , \I0/high/ncd[3] , 
        \I0/high/ncd[2] , \I0/high/ncd[1] , \I0/high/ncd[0] , \I0/high/ba , 
        \I0/high/latch , \I0/high/acb , \I0/high/ctrlack_internal , 
        \I0/high/nlocalcd , \I0/high/U4/U28/U1/clr , \I0/high/U4/U28/U1/set , 
        \I0/high/U1/Z , \I0/high/U1664/y[0] , \I0/high/U1664/y[1] , 
        \I0/high/U1664/x[1] , \I0/high/U1664/x[3] , \I0/high/U1664/x[2] , 
        \I0/high/U1664/x[0] , \I0/high/U1664/U28/Z , \I0/high/U1664/U32/Z , 
        \I0/high/U1664/U29/Z , \I0/high/U1664/U33/Z , \I0/high/U1664/U30/Z , 
        \I0/high/U1664/U31/Z , \I0/high/U1664/U37/Z , \I0/high/U1669/nr , 
        \I0/high/U1669/nd , \I0/high/U1669/n2 , \I1/net20 , \I1/net33 , 
        \I1/net32 , \I1/low/drivel , \I1/low/driveh , \I1/low/localcd , 
        \I1/low/ncd[7] , \I1/low/ncd[6] , \I1/low/ncd[5] , \I1/low/ncd[4] , 
        \I1/low/ncd[3] , \I1/low/ncd[2] , \I1/low/ncd[1] , \I1/low/ncd[0] , 
        \I1/low/ba , \I1/low/latch , \I1/low/acb , \I1/low/ctrlack_internal , 
        \I1/low/nlocalcd , \I1/low/U4/U28/U1/clr , \I1/low/U4/U28/U1/set , 
        \I1/low/U1/Z , \I1/low/U1664/y[0] , \I1/low/U1664/y[1] , 
        \I1/low/U1664/x[1] , \I1/low/U1664/x[3] , \I1/low/U1664/x[2] , 
        \I1/low/U1664/x[0] , \I1/low/U1664/U28/Z , \I1/low/U1664/U32/Z , 
        \I1/low/U1664/U29/Z , \I1/low/U1664/U33/Z , \I1/low/U1664/U30/Z , 
        \I1/low/U1664/U31/Z , \I1/low/U1664/U37/Z , \I1/low/U1669/nr , 
        \I1/low/U1669/nd , \I1/low/U1669/n2 , \I1/high/localcd , 
        \I1/high/ncd[7] , \I1/high/ncd[6] , \I1/high/ncd[5] , \I1/high/ncd[4] , 
        \I1/high/ncd[3] , \I1/high/ncd[2] , \I1/high/ncd[1] , \I1/high/ncd[0] , 
        \I1/high/ba , \I1/high/latch , \I1/high/acb , 
        \I1/high/ctrlack_internal , \I1/high/nlocalcd , 
        \I1/high/U4/U28/U1/clr , \I1/high/U4/U28/U1/set , \I1/high/U1/Z , 
        \I1/high/U1664/y[0] , \I1/high/U1664/y[1] , \I1/high/U1664/x[1] , 
        \I1/high/U1664/x[3] , \I1/high/U1664/x[2] , \I1/high/U1664/x[0] , 
        \I1/high/U1664/U28/Z , \I1/high/U1664/U32/Z , \I1/high/U1664/U29/Z , 
        \I1/high/U1664/U33/Z , \I1/high/U1664/U30/Z , \I1/high/U1664/U31/Z , 
        \I1/high/U1664/U37/Z , \I1/high/U1669/nr , \I1/high/U1669/nd , 
        \I1/high/U1669/n2 , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
    nand2_1 \U3/U5  ( .x(pullreq), .a(net30), .b(net31) );
    nor2_1 \I0/U3/U5  ( .x(net30), .a(\I0/net32 ), .b(\I0/net33 ) );
    buf_2 \I0/low/U1653  ( .x(\I0/low/latch ), .a(\I0/net32 ) );
    nor2_1 \I0/low/U264/U5  ( .x(\I0/low/nlocalcd ), .a(reset), .b(
        \I0/low/localcd ) );
    nor2_1 \I0/low/U1659_0_/U5  ( .x(\I0/low/ncd[0] ), .a(ol[0]), .b(oh[0]) );
    nor2_1 \I0/low/U1659_1_/U5  ( .x(\I0/low/ncd[1] ), .a(ol[1]), .b(oh[1]) );
    nor2_1 \I0/low/U1659_2_/U5  ( .x(\I0/low/ncd[2] ), .a(ol[2]), .b(oh[2]) );
    nor2_1 \I0/low/U1659_3_/U5  ( .x(\I0/low/ncd[3] ), .a(ol[3]), .b(oh[3]) );
    nor2_1 \I0/low/U1659_4_/U5  ( .x(\I0/low/ncd[4] ), .a(ol[4]), .b(oh[4]) );
    nor2_1 \I0/low/U1659_5_/U5  ( .x(\I0/low/ncd[5] ), .a(ol[5]), .b(oh[5]) );
    nor2_1 \I0/low/U1659_6_/U5  ( .x(\I0/low/ncd[6] ), .a(ol[6]), .b(oh[6]) );
    nor2_1 \I0/low/U1659_7_/U5  ( .x(\I0/low/ncd[7] ), .a(ol[7]), .b(oh[7]) );
    nor2_1 \I0/low/U3/U5  ( .x(\I0/low/ctrlack_internal ), .a(\I0/low/acb ), 
        .b(\I0/low/ba ) );
    buf_2 \I0/low/U1665/U7  ( .x(\I0/low/driveh ), .a(\I0/net20 ) );
    buf_2 \I0/low/U1666/U7  ( .x(\I0/low/drivel ), .a(\I0/net20 ) );
    ao23_1 \I0/low/U1658_0_/U21/U1/U1  ( .x(ol[0]), .a(\I0/low/driveh ), .b(ol
        [0]), .c(n1), .d(pull_l[0]), .e(n2) );
    ao23_1 \I0/low/U1658_1_/U21/U1/U1  ( .x(ol[1]), .a(\I0/low/drivel ), .b(ol
        [1]), .c(\I0/low/driveh ), .d(pull_l[1]), .e(n2) );
    ao23_1 \I0/low/U1658_2_/U21/U1/U1  ( .x(ol[2]), .a(\I0/low/drivel ), .b(ol
        [2]), .c(\I0/low/driveh ), .d(pull_l[2]), .e(n2) );
    ao23_1 \I0/low/U1658_3_/U21/U1/U1  ( .x(ol[3]), .a(\I0/low/driveh ), .b(ol
        [3]), .c(\I0/low/drivel ), .d(pull_l[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_4_/U21/U1/U1  ( .x(ol[4]), .a(n1), .b(ol[4]), .c(
        \I0/low/drivel ), .d(pull_l[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_5_/U21/U1/U1  ( .x(ol[5]), .a(\I0/low/driveh ), .b(ol
        [5]), .c(n1), .d(pull_l[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_6_/U21/U1/U1  ( .x(ol[6]), .a(\I0/low/drivel ), .b(ol
        [6]), .c(\I0/low/driveh ), .d(pull_l[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_7_/U21/U1/U1  ( .x(ol[7]), .a(n1), .b(ol[7]), .c(n1), 
        .d(pull_l[7]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_0_/U21/U1/U1  ( .x(oh[0]), .a(\I0/low/driveh ), .b(oh
        [0]), .c(n1), .d(pull_h[0]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_1_/U21/U1/U1  ( .x(oh[1]), .a(n1), .b(oh[1]), .c(
        \I0/low/drivel ), .d(pull_h[1]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_2_/U21/U1/U1  ( .x(oh[2]), .a(\I0/low/drivel ), .b(oh
        [2]), .c(\I0/low/drivel ), .d(pull_h[2]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_3_/U21/U1/U1  ( .x(oh[3]), .a(n1), .b(oh[3]), .c(
        \I0/low/driveh ), .d(pull_h[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_4_/U21/U1/U1  ( .x(oh[4]), .a(n1), .b(oh[4]), .c(n1), 
        .d(pull_h[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_5_/U21/U1/U1  ( .x(oh[5]), .a(\I0/low/drivel ), .b(oh
        [5]), .c(n1), .d(pull_h[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_6_/U21/U1/U1  ( .x(oh[6]), .a(\I0/low/drivel ), .b(oh
        [6]), .c(\I0/low/driveh ), .d(pull_h[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_7_/U21/U1/U1  ( .x(oh[7]), .a(\I0/low/driveh ), .b(oh
        [7]), .c(\I0/low/drivel ), .d(pull_h[7]), .e(\I0/low/latch ) );
    aoai211_1 \I0/low/U4/U28/U1/U1  ( .x(\I0/low/U4/U28/U1/clr ), .a(
        \I0/net20 ), .b(\I0/low/acb ), .c(\I0/low/nlocalcd ), .d(\I0/net32 )
         );
    nand3_1 \I0/low/U4/U28/U1/U2  ( .x(\I0/low/U4/U28/U1/set ), .a(
        \I0/low/nlocalcd ), .b(\I0/net20 ), .c(\I0/low/acb ) );
    nand2_2 \I0/low/U4/U28/U1/U3  ( .x(\I0/net32 ), .a(\I0/low/U4/U28/U1/clr ), 
        .b(\I0/low/U4/U28/U1/set ) );
    oai21_1 \I0/low/U1/U30/U1/U1  ( .x(\I0/low/acb ), .a(\I0/low/U1/Z ), .b(
        \I0/low/ba ), .c(\I0/net20 ) );
    inv_1 \I0/low/U1/U30/U1/U2  ( .x(\I0/low/U1/Z ), .a(\I0/low/acb ) );
    ao222_1 \I0/low/U5/U18/U1/U1  ( .x(\I0/low/ba ), .a(\I0/low/latch ), .b(
        pullcd), .c(\I0/low/latch ), .d(\I0/low/ba ), .e(pullcd), .f(
        \I0/low/ba ) );
    aoi222_1 \I0/low/U1664/U28/U30/U1  ( .x(\I0/low/U1664/x[3] ), .a(
        \I0/low/ncd[7] ), .b(\I0/low/ncd[6] ), .c(\I0/low/ncd[7] ), .d(
        \I0/low/U1664/U28/Z ), .e(\I0/low/ncd[6] ), .f(\I0/low/U1664/U28/Z )
         );
    inv_1 \I0/low/U1664/U28/U30/Uinv  ( .x(\I0/low/U1664/U28/Z ), .a(
        \I0/low/U1664/x[3] ) );
    aoi222_1 \I0/low/U1664/U32/U30/U1  ( .x(\I0/low/U1664/x[0] ), .a(
        \I0/low/ncd[1] ), .b(\I0/low/ncd[0] ), .c(\I0/low/ncd[1] ), .d(
        \I0/low/U1664/U32/Z ), .e(\I0/low/ncd[0] ), .f(\I0/low/U1664/U32/Z )
         );
    inv_1 \I0/low/U1664/U32/U30/Uinv  ( .x(\I0/low/U1664/U32/Z ), .a(
        \I0/low/U1664/x[0] ) );
    aoi222_1 \I0/low/U1664/U29/U30/U1  ( .x(\I0/low/U1664/x[2] ), .a(
        \I0/low/ncd[5] ), .b(\I0/low/ncd[4] ), .c(\I0/low/ncd[5] ), .d(
        \I0/low/U1664/U29/Z ), .e(\I0/low/ncd[4] ), .f(\I0/low/U1664/U29/Z )
         );
    inv_1 \I0/low/U1664/U29/U30/Uinv  ( .x(\I0/low/U1664/U29/Z ), .a(
        \I0/low/U1664/x[2] ) );
    aoi222_1 \I0/low/U1664/U33/U30/U1  ( .x(\I0/low/U1664/y[0] ), .a(
        \I0/low/U1664/x[1] ), .b(\I0/low/U1664/x[0] ), .c(\I0/low/U1664/x[1] ), 
        .d(\I0/low/U1664/U33/Z ), .e(\I0/low/U1664/x[0] ), .f(
        \I0/low/U1664/U33/Z ) );
    inv_1 \I0/low/U1664/U33/U30/Uinv  ( .x(\I0/low/U1664/U33/Z ), .a(
        \I0/low/U1664/y[0] ) );
    aoi222_1 \I0/low/U1664/U30/U30/U1  ( .x(\I0/low/U1664/y[1] ), .a(
        \I0/low/U1664/x[3] ), .b(\I0/low/U1664/x[2] ), .c(\I0/low/U1664/x[3] ), 
        .d(\I0/low/U1664/U30/Z ), .e(\I0/low/U1664/x[2] ), .f(
        \I0/low/U1664/U30/Z ) );
    inv_1 \I0/low/U1664/U30/U30/Uinv  ( .x(\I0/low/U1664/U30/Z ), .a(
        \I0/low/U1664/y[1] ) );
    aoi222_1 \I0/low/U1664/U31/U30/U1  ( .x(\I0/low/U1664/x[1] ), .a(
        \I0/low/ncd[3] ), .b(\I0/low/ncd[2] ), .c(\I0/low/ncd[3] ), .d(
        \I0/low/U1664/U31/Z ), .e(\I0/low/ncd[2] ), .f(\I0/low/U1664/U31/Z )
         );
    inv_1 \I0/low/U1664/U31/U30/Uinv  ( .x(\I0/low/U1664/U31/Z ), .a(
        \I0/low/U1664/x[1] ) );
    aoi222_1 \I0/low/U1664/U37/U30/U1  ( .x(\I0/low/localcd ), .a(
        \I0/low/U1664/y[0] ), .b(\I0/low/U1664/y[1] ), .c(\I0/low/U1664/y[0] ), 
        .d(\I0/low/U1664/U37/Z ), .e(\I0/low/U1664/y[1] ), .f(
        \I0/low/U1664/U37/Z ) );
    inv_1 \I0/low/U1664/U37/U30/Uinv  ( .x(\I0/low/U1664/U37/Z ), .a(
        \I0/low/localcd ) );
    nor3_1 \I0/low/U1669/Unr  ( .x(\I0/low/U1669/nr ), .a(
        \I0/low/ctrlack_internal ), .b(n1), .c(\I0/low/driveh ) );
    nand3_1 \I0/low/U1669/Und  ( .x(\I0/low/U1669/nd ), .a(
        \I0/low/ctrlack_internal ), .b(\I0/low/drivel ), .c(\I0/low/driveh )
         );
    oa21_1 \I0/low/U1669/U1  ( .x(\I0/low/U1669/n2 ), .a(\I0/low/U1669/n2 ), 
        .b(\I0/low/U1669/nr ), .c(\I0/low/U1669/nd ) );
    inv_2 \I0/low/U1669/U3  ( .x(ctrlack), .a(\I0/low/U1669/n2 ) );
    buf_2 \I0/high/U1653  ( .x(\I0/high/latch ), .a(\I0/net33 ) );
    nor2_1 \I0/high/U264/U5  ( .x(\I0/high/nlocalcd ), .a(reset), .b(
        \I0/high/localcd ) );
    nor2_1 \I0/high/U1659_0_/U5  ( .x(\I0/high/ncd[0] ), .a(ol[8]), .b(oh[8])
         );
    nor2_1 \I0/high/U1659_1_/U5  ( .x(\I0/high/ncd[1] ), .a(ol[9]), .b(oh[9])
         );
    nor2_1 \I0/high/U1659_2_/U5  ( .x(\I0/high/ncd[2] ), .a(ol[10]), .b(oh[10]
        ) );
    nor2_1 \I0/high/U1659_3_/U5  ( .x(\I0/high/ncd[3] ), .a(ol[11]), .b(oh[11]
        ) );
    nor2_1 \I0/high/U1659_4_/U5  ( .x(\I0/high/ncd[4] ), .a(ol[12]), .b(oh[12]
        ) );
    nor2_1 \I0/high/U1659_5_/U5  ( .x(\I0/high/ncd[5] ), .a(ol[13]), .b(oh[13]
        ) );
    nor2_1 \I0/high/U1659_6_/U5  ( .x(\I0/high/ncd[6] ), .a(ol[14]), .b(oh[14]
        ) );
    nor2_1 \I0/high/U1659_7_/U5  ( .x(\I0/high/ncd[7] ), .a(ol[15]), .b(oh[15]
        ) );
    nor2_1 \I0/high/U3/U5  ( .x(\I0/high/ctrlack_internal ), .a(\I0/high/acb ), 
        .b(\I0/high/ba ) );
    buf_2 \I0/high/U1665/U7  ( .x(\I0/high/driveh ), .a(net17) );
    buf_2 \I0/high/U1666/U7  ( .x(\I0/high/drivel ), .a(net17) );
    ao23_1 \I0/high/U1658_0_/U21/U1/U1  ( .x(ol[8]), .a(\I0/high/driveh ), .b(
        ol[8]), .c(n3), .d(pull_l[0]), .e(n4) );
    ao23_1 \I0/high/U1658_1_/U21/U1/U1  ( .x(ol[9]), .a(\I0/high/drivel ), .b(
        ol[9]), .c(\I0/high/driveh ), .d(pull_l[1]), .e(n4) );
    ao23_1 \I0/high/U1658_2_/U21/U1/U1  ( .x(ol[10]), .a(\I0/high/drivel ), 
        .b(ol[10]), .c(\I0/high/driveh ), .d(pull_l[2]), .e(n4) );
    ao23_1 \I0/high/U1658_3_/U21/U1/U1  ( .x(ol[11]), .a(\I0/high/driveh ), 
        .b(ol[11]), .c(\I0/high/drivel ), .d(pull_l[3]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_4_/U21/U1/U1  ( .x(ol[12]), .a(n3), .b(ol[12]), .c(
        \I0/high/drivel ), .d(pull_l[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_5_/U21/U1/U1  ( .x(ol[13]), .a(\I0/high/driveh ), 
        .b(ol[13]), .c(n3), .d(pull_l[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_6_/U21/U1/U1  ( .x(ol[14]), .a(\I0/high/drivel ), 
        .b(ol[14]), .c(\I0/high/driveh ), .d(pull_l[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_7_/U21/U1/U1  ( .x(ol[15]), .a(n3), .b(ol[15]), .c(
        n3), .d(pull_l[7]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_0_/U21/U1/U1  ( .x(oh[8]), .a(\I0/high/driveh ), .b(
        oh[8]), .c(n3), .d(pull_h[0]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_1_/U21/U1/U1  ( .x(oh[9]), .a(n3), .b(oh[9]), .c(
        \I0/high/drivel ), .d(pull_h[1]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_2_/U21/U1/U1  ( .x(oh[10]), .a(\I0/high/drivel ), 
        .b(oh[10]), .c(\I0/high/drivel ), .d(pull_h[2]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_3_/U21/U1/U1  ( .x(oh[11]), .a(n3), .b(oh[11]), .c(
        \I0/high/driveh ), .d(pull_h[3]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_4_/U21/U1/U1  ( .x(oh[12]), .a(n3), .b(oh[12]), .c(
        n3), .d(pull_h[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_5_/U21/U1/U1  ( .x(oh[13]), .a(\I0/high/drivel ), 
        .b(oh[13]), .c(n3), .d(pull_h[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_6_/U21/U1/U1  ( .x(oh[14]), .a(\I0/high/drivel ), 
        .b(oh[14]), .c(\I0/high/driveh ), .d(pull_h[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_7_/U21/U1/U1  ( .x(oh[15]), .a(\I0/high/driveh ), 
        .b(oh[15]), .c(\I0/high/drivel ), .d(pull_h[7]), .e(\I0/high/latch )
         );
    aoai211_1 \I0/high/U4/U28/U1/U1  ( .x(\I0/high/U4/U28/U1/clr ), .a(net17), 
        .b(\I0/high/acb ), .c(\I0/high/nlocalcd ), .d(\I0/net33 ) );
    nand3_1 \I0/high/U4/U28/U1/U2  ( .x(\I0/high/U4/U28/U1/set ), .a(
        \I0/high/nlocalcd ), .b(net17), .c(\I0/high/acb ) );
    nand2_2 \I0/high/U4/U28/U1/U3  ( .x(\I0/net33 ), .a(
        \I0/high/U4/U28/U1/clr ), .b(\I0/high/U4/U28/U1/set ) );
    oai21_1 \I0/high/U1/U30/U1/U1  ( .x(\I0/high/acb ), .a(\I0/high/U1/Z ), 
        .b(\I0/high/ba ), .c(net17) );
    inv_1 \I0/high/U1/U30/U1/U2  ( .x(\I0/high/U1/Z ), .a(\I0/high/acb ) );
    ao222_1 \I0/high/U5/U18/U1/U1  ( .x(\I0/high/ba ), .a(\I0/high/latch ), 
        .b(pullcd), .c(\I0/high/latch ), .d(\I0/high/ba ), .e(pullcd), .f(
        \I0/high/ba ) );
    aoi222_1 \I0/high/U1664/U28/U30/U1  ( .x(\I0/high/U1664/x[3] ), .a(
        \I0/high/ncd[7] ), .b(\I0/high/ncd[6] ), .c(\I0/high/ncd[7] ), .d(
        \I0/high/U1664/U28/Z ), .e(\I0/high/ncd[6] ), .f(\I0/high/U1664/U28/Z 
        ) );
    inv_1 \I0/high/U1664/U28/U30/Uinv  ( .x(\I0/high/U1664/U28/Z ), .a(
        \I0/high/U1664/x[3] ) );
    aoi222_1 \I0/high/U1664/U32/U30/U1  ( .x(\I0/high/U1664/x[0] ), .a(
        \I0/high/ncd[1] ), .b(\I0/high/ncd[0] ), .c(\I0/high/ncd[1] ), .d(
        \I0/high/U1664/U32/Z ), .e(\I0/high/ncd[0] ), .f(\I0/high/U1664/U32/Z 
        ) );
    inv_1 \I0/high/U1664/U32/U30/Uinv  ( .x(\I0/high/U1664/U32/Z ), .a(
        \I0/high/U1664/x[0] ) );
    aoi222_1 \I0/high/U1664/U29/U30/U1  ( .x(\I0/high/U1664/x[2] ), .a(
        \I0/high/ncd[5] ), .b(\I0/high/ncd[4] ), .c(\I0/high/ncd[5] ), .d(
        \I0/high/U1664/U29/Z ), .e(\I0/high/ncd[4] ), .f(\I0/high/U1664/U29/Z 
        ) );
    inv_1 \I0/high/U1664/U29/U30/Uinv  ( .x(\I0/high/U1664/U29/Z ), .a(
        \I0/high/U1664/x[2] ) );
    aoi222_1 \I0/high/U1664/U33/U30/U1  ( .x(\I0/high/U1664/y[0] ), .a(
        \I0/high/U1664/x[1] ), .b(\I0/high/U1664/x[0] ), .c(
        \I0/high/U1664/x[1] ), .d(\I0/high/U1664/U33/Z ), .e(
        \I0/high/U1664/x[0] ), .f(\I0/high/U1664/U33/Z ) );
    inv_1 \I0/high/U1664/U33/U30/Uinv  ( .x(\I0/high/U1664/U33/Z ), .a(
        \I0/high/U1664/y[0] ) );
    aoi222_1 \I0/high/U1664/U30/U30/U1  ( .x(\I0/high/U1664/y[1] ), .a(
        \I0/high/U1664/x[3] ), .b(\I0/high/U1664/x[2] ), .c(
        \I0/high/U1664/x[3] ), .d(\I0/high/U1664/U30/Z ), .e(
        \I0/high/U1664/x[2] ), .f(\I0/high/U1664/U30/Z ) );
    inv_1 \I0/high/U1664/U30/U30/Uinv  ( .x(\I0/high/U1664/U30/Z ), .a(
        \I0/high/U1664/y[1] ) );
    aoi222_1 \I0/high/U1664/U31/U30/U1  ( .x(\I0/high/U1664/x[1] ), .a(
        \I0/high/ncd[3] ), .b(\I0/high/ncd[2] ), .c(\I0/high/ncd[3] ), .d(
        \I0/high/U1664/U31/Z ), .e(\I0/high/ncd[2] ), .f(\I0/high/U1664/U31/Z 
        ) );
    inv_1 \I0/high/U1664/U31/U30/Uinv  ( .x(\I0/high/U1664/U31/Z ), .a(
        \I0/high/U1664/x[1] ) );
    aoi222_1 \I0/high/U1664/U37/U30/U1  ( .x(\I0/high/localcd ), .a(
        \I0/high/U1664/y[0] ), .b(\I0/high/U1664/y[1] ), .c(
        \I0/high/U1664/y[0] ), .d(\I0/high/U1664/U37/Z ), .e(
        \I0/high/U1664/y[1] ), .f(\I0/high/U1664/U37/Z ) );
    inv_1 \I0/high/U1664/U37/U30/Uinv  ( .x(\I0/high/U1664/U37/Z ), .a(
        \I0/high/localcd ) );
    nor3_1 \I0/high/U1669/Unr  ( .x(\I0/high/U1669/nr ), .a(
        \I0/high/ctrlack_internal ), .b(n3), .c(\I0/high/driveh ) );
    nand3_1 \I0/high/U1669/Und  ( .x(\I0/high/U1669/nd ), .a(
        \I0/high/ctrlack_internal ), .b(\I0/high/drivel ), .c(\I0/high/driveh 
        ) );
    oa21_1 \I0/high/U1669/U1  ( .x(\I0/high/U1669/n2 ), .a(\I0/high/U1669/n2 ), 
        .b(\I0/high/U1669/nr ), .c(\I0/high/U1669/nd ) );
    inv_2 \I0/high/U1669/U3  ( .x(\I0/net20 ), .a(\I0/high/U1669/n2 ) );
    nor2_1 \I1/U3/U5  ( .x(net31), .a(\I1/net32 ), .b(\I1/net33 ) );
    buf_2 \I1/low/U1653  ( .x(\I1/low/latch ), .a(\I1/net32 ) );
    nor2_1 \I1/low/U264/U5  ( .x(\I1/low/nlocalcd ), .a(reset), .b(
        \I1/low/localcd ) );
    nor2_1 \I1/low/U1659_0_/U5  ( .x(\I1/low/ncd[0] ), .a(ol[16]), .b(oh[16])
         );
    nor2_1 \I1/low/U1659_1_/U5  ( .x(\I1/low/ncd[1] ), .a(ol[17]), .b(oh[17])
         );
    nor2_1 \I1/low/U1659_2_/U5  ( .x(\I1/low/ncd[2] ), .a(ol[18]), .b(oh[18])
         );
    nor2_1 \I1/low/U1659_3_/U5  ( .x(\I1/low/ncd[3] ), .a(ol[19]), .b(oh[19])
         );
    nor2_1 \I1/low/U1659_4_/U5  ( .x(\I1/low/ncd[4] ), .a(ol[20]), .b(oh[20])
         );
    nor2_1 \I1/low/U1659_5_/U5  ( .x(\I1/low/ncd[5] ), .a(ol[21]), .b(oh[21])
         );
    nor2_1 \I1/low/U1659_6_/U5  ( .x(\I1/low/ncd[6] ), .a(ol[22]), .b(oh[22])
         );
    nor2_1 \I1/low/U1659_7_/U5  ( .x(\I1/low/ncd[7] ), .a(ol[23]), .b(oh[23])
         );
    nor2_1 \I1/low/U3/U5  ( .x(\I1/low/ctrlack_internal ), .a(\I1/low/acb ), 
        .b(\I1/low/ba ) );
    buf_2 \I1/low/U1665/U7  ( .x(\I1/low/driveh ), .a(\I1/net20 ) );
    buf_2 \I1/low/U1666/U7  ( .x(\I1/low/drivel ), .a(\I1/net20 ) );
    ao23_1 \I1/low/U1658_0_/U21/U1/U1  ( .x(ol[16]), .a(\I1/low/drivel ), .b(
        ol[16]), .c(n5), .d(pull_l[0]), .e(n6) );
    ao23_1 \I1/low/U1658_1_/U21/U1/U1  ( .x(ol[17]), .a(\I1/low/driveh ), .b(
        ol[17]), .c(n5), .d(pull_l[1]), .e(n6) );
    ao23_1 \I1/low/U1658_2_/U21/U1/U1  ( .x(ol[18]), .a(\I1/low/drivel ), .b(
        ol[18]), .c(\I1/low/driveh ), .d(pull_l[2]), .e(n6) );
    ao23_1 \I1/low/U1658_3_/U21/U1/U1  ( .x(ol[19]), .a(n5), .b(ol[19]), .c(
        \I1/low/driveh ), .d(pull_l[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_4_/U21/U1/U1  ( .x(ol[20]), .a(\I1/low/driveh ), .b(
        ol[20]), .c(\I1/low/drivel ), .d(pull_l[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_5_/U21/U1/U1  ( .x(ol[21]), .a(n5), .b(ol[21]), .c(
        \I1/low/drivel ), .d(pull_l[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_6_/U21/U1/U1  ( .x(ol[22]), .a(\I1/low/driveh ), .b(
        ol[22]), .c(n5), .d(pull_l[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_7_/U21/U1/U1  ( .x(ol[23]), .a(\I1/low/drivel ), .b(
        ol[23]), .c(\I1/low/driveh ), .d(pull_l[7]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_0_/U21/U1/U1  ( .x(oh[16]), .a(\I1/low/driveh ), .b(
        oh[16]), .c(\I1/low/drivel ), .d(pull_h[0]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_1_/U21/U1/U1  ( .x(oh[17]), .a(\I1/low/drivel ), .b(
        oh[17]), .c(n5), .d(pull_h[1]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_2_/U21/U1/U1  ( .x(oh[18]), .a(\I1/low/drivel ), .b(
        oh[18]), .c(\I1/low/driveh ), .d(pull_h[2]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_3_/U21/U1/U1  ( .x(oh[19]), .a(n5), .b(oh[19]), .c(n5
        ), .d(pull_h[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_4_/U21/U1/U1  ( .x(oh[20]), .a(n5), .b(oh[20]), .c(n5
        ), .d(pull_h[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_5_/U21/U1/U1  ( .x(oh[21]), .a(\I1/low/drivel ), .b(
        oh[21]), .c(\I1/low/driveh ), .d(pull_h[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_6_/U21/U1/U1  ( .x(oh[22]), .a(n5), .b(oh[22]), .c(
        \I1/low/drivel ), .d(pull_h[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_7_/U21/U1/U1  ( .x(oh[23]), .a(\I1/low/driveh ), .b(
        oh[23]), .c(\I1/low/drivel ), .d(pull_h[7]), .e(\I1/low/latch ) );
    aoai211_1 \I1/low/U4/U28/U1/U1  ( .x(\I1/low/U4/U28/U1/clr ), .a(
        \I1/net20 ), .b(\I1/low/acb ), .c(\I1/low/nlocalcd ), .d(\I1/net32 )
         );
    nand3_1 \I1/low/U4/U28/U1/U2  ( .x(\I1/low/U4/U28/U1/set ), .a(
        \I1/low/nlocalcd ), .b(\I1/net20 ), .c(\I1/low/acb ) );
    nand2_2 \I1/low/U4/U28/U1/U3  ( .x(\I1/net32 ), .a(\I1/low/U4/U28/U1/clr ), 
        .b(\I1/low/U4/U28/U1/set ) );
    oai21_1 \I1/low/U1/U30/U1/U1  ( .x(\I1/low/acb ), .a(\I1/low/U1/Z ), .b(
        \I1/low/ba ), .c(\I1/net20 ) );
    inv_1 \I1/low/U1/U30/U1/U2  ( .x(\I1/low/U1/Z ), .a(\I1/low/acb ) );
    ao222_1 \I1/low/U5/U18/U1/U1  ( .x(\I1/low/ba ), .a(\I1/low/latch ), .b(
        pullcd), .c(\I1/low/latch ), .d(\I1/low/ba ), .e(pullcd), .f(
        \I1/low/ba ) );
    aoi222_1 \I1/low/U1664/U28/U30/U1  ( .x(\I1/low/U1664/x[3] ), .a(
        \I1/low/ncd[7] ), .b(\I1/low/ncd[6] ), .c(\I1/low/ncd[7] ), .d(
        \I1/low/U1664/U28/Z ), .e(\I1/low/ncd[6] ), .f(\I1/low/U1664/U28/Z )
         );
    inv_1 \I1/low/U1664/U28/U30/Uinv  ( .x(\I1/low/U1664/U28/Z ), .a(
        \I1/low/U1664/x[3] ) );
    aoi222_1 \I1/low/U1664/U32/U30/U1  ( .x(\I1/low/U1664/x[0] ), .a(
        \I1/low/ncd[1] ), .b(\I1/low/ncd[0] ), .c(\I1/low/ncd[1] ), .d(
        \I1/low/U1664/U32/Z ), .e(\I1/low/ncd[0] ), .f(\I1/low/U1664/U32/Z )
         );
    inv_1 \I1/low/U1664/U32/U30/Uinv  ( .x(\I1/low/U1664/U32/Z ), .a(
        \I1/low/U1664/x[0] ) );
    aoi222_1 \I1/low/U1664/U29/U30/U1  ( .x(\I1/low/U1664/x[2] ), .a(
        \I1/low/ncd[5] ), .b(\I1/low/ncd[4] ), .c(\I1/low/ncd[5] ), .d(
        \I1/low/U1664/U29/Z ), .e(\I1/low/ncd[4] ), .f(\I1/low/U1664/U29/Z )
         );
    inv_1 \I1/low/U1664/U29/U30/Uinv  ( .x(\I1/low/U1664/U29/Z ), .a(
        \I1/low/U1664/x[2] ) );
    aoi222_1 \I1/low/U1664/U33/U30/U1  ( .x(\I1/low/U1664/y[0] ), .a(
        \I1/low/U1664/x[1] ), .b(\I1/low/U1664/x[0] ), .c(\I1/low/U1664/x[1] ), 
        .d(\I1/low/U1664/U33/Z ), .e(\I1/low/U1664/x[0] ), .f(
        \I1/low/U1664/U33/Z ) );
    inv_1 \I1/low/U1664/U33/U30/Uinv  ( .x(\I1/low/U1664/U33/Z ), .a(
        \I1/low/U1664/y[0] ) );
    aoi222_1 \I1/low/U1664/U30/U30/U1  ( .x(\I1/low/U1664/y[1] ), .a(
        \I1/low/U1664/x[3] ), .b(\I1/low/U1664/x[2] ), .c(\I1/low/U1664/x[3] ), 
        .d(\I1/low/U1664/U30/Z ), .e(\I1/low/U1664/x[2] ), .f(
        \I1/low/U1664/U30/Z ) );
    inv_1 \I1/low/U1664/U30/U30/Uinv  ( .x(\I1/low/U1664/U30/Z ), .a(
        \I1/low/U1664/y[1] ) );
    aoi222_1 \I1/low/U1664/U31/U30/U1  ( .x(\I1/low/U1664/x[1] ), .a(
        \I1/low/ncd[3] ), .b(\I1/low/ncd[2] ), .c(\I1/low/ncd[3] ), .d(
        \I1/low/U1664/U31/Z ), .e(\I1/low/ncd[2] ), .f(\I1/low/U1664/U31/Z )
         );
    inv_1 \I1/low/U1664/U31/U30/Uinv  ( .x(\I1/low/U1664/U31/Z ), .a(
        \I1/low/U1664/x[1] ) );
    aoi222_1 \I1/low/U1664/U37/U30/U1  ( .x(\I1/low/localcd ), .a(
        \I1/low/U1664/y[0] ), .b(\I1/low/U1664/y[1] ), .c(\I1/low/U1664/y[0] ), 
        .d(\I1/low/U1664/U37/Z ), .e(\I1/low/U1664/y[1] ), .f(
        \I1/low/U1664/U37/Z ) );
    inv_1 \I1/low/U1664/U37/U30/Uinv  ( .x(\I1/low/U1664/U37/Z ), .a(
        \I1/low/localcd ) );
    nor3_1 \I1/low/U1669/Unr  ( .x(\I1/low/U1669/nr ), .a(
        \I1/low/ctrlack_internal ), .b(n5), .c(\I1/low/driveh ) );
    nand3_1 \I1/low/U1669/Und  ( .x(\I1/low/U1669/nd ), .a(
        \I1/low/ctrlack_internal ), .b(\I1/low/drivel ), .c(\I1/low/driveh )
         );
    oa21_1 \I1/low/U1669/U1  ( .x(\I1/low/U1669/n2 ), .a(\I1/low/U1669/n2 ), 
        .b(\I1/low/U1669/nr ), .c(\I1/low/U1669/nd ) );
    inv_2 \I1/low/U1669/U3  ( .x(net17), .a(\I1/low/U1669/n2 ) );
    buf_2 \I1/high/U1653  ( .x(\I1/high/latch ), .a(\I1/net33 ) );
    nor2_1 \I1/high/U264/U5  ( .x(\I1/high/nlocalcd ), .a(reset), .b(
        \I1/high/localcd ) );
    nor2_1 \I1/high/U1659_0_/U5  ( .x(\I1/high/ncd[0] ), .a(ol[24]), .b(oh[24]
        ) );
    nor2_1 \I1/high/U1659_1_/U5  ( .x(\I1/high/ncd[1] ), .a(ol[25]), .b(oh[25]
        ) );
    nor2_1 \I1/high/U1659_2_/U5  ( .x(\I1/high/ncd[2] ), .a(ol[26]), .b(oh[26]
        ) );
    nor2_1 \I1/high/U1659_3_/U5  ( .x(\I1/high/ncd[3] ), .a(ol[27]), .b(oh[27]
        ) );
    nor2_1 \I1/high/U1659_4_/U5  ( .x(\I1/high/ncd[4] ), .a(ol[28]), .b(oh[28]
        ) );
    nor2_1 \I1/high/U1659_5_/U5  ( .x(\I1/high/ncd[5] ), .a(ol[29]), .b(oh[29]
        ) );
    nor2_1 \I1/high/U1659_6_/U5  ( .x(\I1/high/ncd[6] ), .a(ol[30]), .b(oh[30]
        ) );
    nor2_1 \I1/high/U1659_7_/U5  ( .x(\I1/high/ncd[7] ), .a(ol[31]), .b(oh[31]
        ) );
    nor2_1 \I1/high/U3/U5  ( .x(\I1/high/ctrlack_internal ), .a(\I1/high/acb ), 
        .b(\I1/high/ba ) );
    ao23_1 \I1/high/U1658_0_/U21/U1/U1  ( .x(ol[24]), .a(n7), .b(ol[24]), .c(
        n8), .d(pull_l[0]), .e(n12) );
    ao23_1 \I1/high/U1658_1_/U21/U1/U1  ( .x(ol[25]), .a(n7), .b(ol[25]), .c(
        n8), .d(pull_l[1]), .e(n12) );
    ao23_1 \I1/high/U1658_2_/U21/U1/U1  ( .x(ol[26]), .a(n7), .b(ol[26]), .c(
        n7), .d(pull_l[2]), .e(n12) );
    ao23_1 \I1/high/U1658_3_/U21/U1/U1  ( .x(ol[27]), .a(n7), .b(ol[27]), .c(
        n7), .d(pull_l[3]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_4_/U21/U1/U1  ( .x(ol[28]), .a(n7), .b(ol[28]), .c(
        n7), .d(pull_l[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_5_/U21/U1/U1  ( .x(ol[29]), .a(n7), .b(ol[29]), .c(
        n8), .d(pull_l[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_6_/U21/U1/U1  ( .x(ol[30]), .a(n7), .b(ol[30]), .c(
        n8), .d(pull_l[6]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_7_/U21/U1/U1  ( .x(ol[31]), .a(n7), .b(ol[31]), .c(
        n8), .d(pull_l[7]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_0_/U21/U1/U1  ( .x(oh[24]), .a(n10), .b(oh[24]), .c(
        n10), .d(pull_h[0]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_1_/U21/U1/U1  ( .x(oh[25]), .a(n10), .b(oh[25]), .c(
        n11), .d(pull_h[1]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_2_/U21/U1/U1  ( .x(oh[26]), .a(n10), .b(oh[26]), .c(
        n11), .d(pull_h[2]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_3_/U21/U1/U1  ( .x(oh[27]), .a(n10), .b(oh[27]), .c(
        n10), .d(pull_h[3]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_4_/U21/U1/U1  ( .x(oh[28]), .a(n10), .b(oh[28]), .c(
        n11), .d(pull_h[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_5_/U21/U1/U1  ( .x(oh[29]), .a(n10), .b(oh[29]), .c(
        n11), .d(pull_h[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_6_/U21/U1/U1  ( .x(oh[30]), .a(n10), .b(oh[30]), .c(
        n11), .d(pull_h[6]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_7_/U21/U1/U1  ( .x(oh[31]), .a(n10), .b(oh[31]), .c(
        n10), .d(pull_h[7]), .e(\I1/high/latch ) );
    aoai211_1 \I1/high/U4/U28/U1/U1  ( .x(\I1/high/U4/U28/U1/clr ), .a(ctrlreq
        ), .b(\I1/high/acb ), .c(\I1/high/nlocalcd ), .d(\I1/net33 ) );
    nand3_1 \I1/high/U4/U28/U1/U2  ( .x(\I1/high/U4/U28/U1/set ), .a(
        \I1/high/nlocalcd ), .b(ctrlreq), .c(\I1/high/acb ) );
    nand2_2 \I1/high/U4/U28/U1/U3  ( .x(\I1/net33 ), .a(
        \I1/high/U4/U28/U1/clr ), .b(\I1/high/U4/U28/U1/set ) );
    oai21_1 \I1/high/U1/U30/U1/U1  ( .x(\I1/high/acb ), .a(\I1/high/U1/Z ), 
        .b(\I1/high/ba ), .c(ctrlreq) );
    inv_1 \I1/high/U1/U30/U1/U2  ( .x(\I1/high/U1/Z ), .a(\I1/high/acb ) );
    ao222_1 \I1/high/U5/U18/U1/U1  ( .x(\I1/high/ba ), .a(\I1/high/latch ), 
        .b(pullcd), .c(\I1/high/latch ), .d(\I1/high/ba ), .e(pullcd), .f(
        \I1/high/ba ) );
    aoi222_1 \I1/high/U1664/U28/U30/U1  ( .x(\I1/high/U1664/x[3] ), .a(
        \I1/high/ncd[7] ), .b(\I1/high/ncd[6] ), .c(\I1/high/ncd[7] ), .d(
        \I1/high/U1664/U28/Z ), .e(\I1/high/ncd[6] ), .f(\I1/high/U1664/U28/Z 
        ) );
    inv_1 \I1/high/U1664/U28/U30/Uinv  ( .x(\I1/high/U1664/U28/Z ), .a(
        \I1/high/U1664/x[3] ) );
    aoi222_1 \I1/high/U1664/U32/U30/U1  ( .x(\I1/high/U1664/x[0] ), .a(
        \I1/high/ncd[1] ), .b(\I1/high/ncd[0] ), .c(\I1/high/ncd[1] ), .d(
        \I1/high/U1664/U32/Z ), .e(\I1/high/ncd[0] ), .f(\I1/high/U1664/U32/Z 
        ) );
    inv_1 \I1/high/U1664/U32/U30/Uinv  ( .x(\I1/high/U1664/U32/Z ), .a(
        \I1/high/U1664/x[0] ) );
    aoi222_1 \I1/high/U1664/U29/U30/U1  ( .x(\I1/high/U1664/x[2] ), .a(
        \I1/high/ncd[5] ), .b(\I1/high/ncd[4] ), .c(\I1/high/ncd[5] ), .d(
        \I1/high/U1664/U29/Z ), .e(\I1/high/ncd[4] ), .f(\I1/high/U1664/U29/Z 
        ) );
    inv_1 \I1/high/U1664/U29/U30/Uinv  ( .x(\I1/high/U1664/U29/Z ), .a(
        \I1/high/U1664/x[2] ) );
    aoi222_1 \I1/high/U1664/U33/U30/U1  ( .x(\I1/high/U1664/y[0] ), .a(
        \I1/high/U1664/x[1] ), .b(\I1/high/U1664/x[0] ), .c(
        \I1/high/U1664/x[1] ), .d(\I1/high/U1664/U33/Z ), .e(
        \I1/high/U1664/x[0] ), .f(\I1/high/U1664/U33/Z ) );
    inv_1 \I1/high/U1664/U33/U30/Uinv  ( .x(\I1/high/U1664/U33/Z ), .a(
        \I1/high/U1664/y[0] ) );
    aoi222_1 \I1/high/U1664/U30/U30/U1  ( .x(\I1/high/U1664/y[1] ), .a(
        \I1/high/U1664/x[3] ), .b(\I1/high/U1664/x[2] ), .c(
        \I1/high/U1664/x[3] ), .d(\I1/high/U1664/U30/Z ), .e(
        \I1/high/U1664/x[2] ), .f(\I1/high/U1664/U30/Z ) );
    inv_1 \I1/high/U1664/U30/U30/Uinv  ( .x(\I1/high/U1664/U30/Z ), .a(
        \I1/high/U1664/y[1] ) );
    aoi222_1 \I1/high/U1664/U31/U30/U1  ( .x(\I1/high/U1664/x[1] ), .a(
        \I1/high/ncd[3] ), .b(\I1/high/ncd[2] ), .c(\I1/high/ncd[3] ), .d(
        \I1/high/U1664/U31/Z ), .e(\I1/high/ncd[2] ), .f(\I1/high/U1664/U31/Z 
        ) );
    inv_1 \I1/high/U1664/U31/U30/Uinv  ( .x(\I1/high/U1664/U31/Z ), .a(
        \I1/high/U1664/x[1] ) );
    aoi222_1 \I1/high/U1664/U37/U30/U1  ( .x(\I1/high/localcd ), .a(
        \I1/high/U1664/y[0] ), .b(\I1/high/U1664/y[1] ), .c(
        \I1/high/U1664/y[0] ), .d(\I1/high/U1664/U37/Z ), .e(
        \I1/high/U1664/y[1] ), .f(\I1/high/U1664/U37/Z ) );
    inv_1 \I1/high/U1664/U37/U30/Uinv  ( .x(\I1/high/U1664/U37/Z ), .a(
        \I1/high/localcd ) );
    nor3_1 \I1/high/U1669/Unr  ( .x(\I1/high/U1669/nr ), .a(
        \I1/high/ctrlack_internal ), .b(n8), .c(n11) );
    nand3_1 \I1/high/U1669/Und  ( .x(\I1/high/U1669/nd ), .a(
        \I1/high/ctrlack_internal ), .b(n8), .c(n11) );
    oa21_1 \I1/high/U1669/U1  ( .x(\I1/high/U1669/n2 ), .a(\I1/high/U1669/n2 ), 
        .b(\I1/high/U1669/nr ), .c(\I1/high/U1669/nd ) );
    inv_2 \I1/high/U1669/U3  ( .x(\I1/net20 ), .a(\I1/high/U1669/n2 ) );
    buf_2 U1 ( .x(n1), .a(\I0/net20 ) );
    buf_1 U2 ( .x(n2), .a(\I0/low/latch ) );
    buf_2 U3 ( .x(n3), .a(net17) );
    buf_1 U4 ( .x(n4), .a(\I0/high/latch ) );
    buf_2 U5 ( .x(n5), .a(\I1/net20 ) );
    buf_1 U6 ( .x(n6), .a(\I1/low/latch ) );
    inv_2 U7 ( .x(n7), .a(n9) );
    inv_1 U8 ( .x(n8), .a(n9) );
    inv_0 U9 ( .x(n9), .a(ctrlreq) );
    inv_2 U10 ( .x(n10), .a(n9) );
    inv_1 U11 ( .x(n11), .a(n9) );
    buf_1 U12 ( .x(n12), .a(\I1/high/latch ) );
endmodule


module chain_fr2dr_byte_2 ( nia, oh, ol, i, nReset, noa );
output [7:0] oh;
output [7:0] ol;
input  [4:0] i;
input  nReset, noa;
output nia;
    wire eop, net135, nca, nbReset, ncla, \c[3] , \c[2] , \c[1] , \c[0] , 
        \cl[3] , \cl[2] , \cl[1] , \cl[0] , asel, bsel, asela, bsela, csel, 
        dsel, csela, dsela, esel, fsel, esela, fsela, naa, nda, \a[3] , \a[2] , 
        \a[1] , \a[0] , \d[3] , \d[2] , \d[1] , \d[0] , nba, nea, nfa, \b[3] , 
        \b[2] , \b[1] , \b[0] , \f[3] , \f[2] , \f[1] , \f[0] , \e[3] , \e[2] , 
        \e[1] , \e[0] , \U891/nack , \U891/acka , \U891/naack[0] , 
        \U891/naack[1] , \U891/iay , \U891/ackb , \U891/reset , \U891/neopack , 
        \U891/U1128/nb , \U891/U1128/na , \U891/U1118_0_/nr , 
        \U891/U1118_0_/nd , \U891/U1118_0_/n2 , \U891/U1118_1_/nr , 
        \U891/U1118_1_/nd , \U891/U1118_1_/n2 , \U891/U1118_2_/nr , 
        \U891/U1118_2_/nd , \U891/U1118_2_/n2 , \U891/U1118_3_/nr , 
        \U891/U1118_3_/nd , \U891/U1118_3_/n2 , \U891/U1117_0_/nr , 
        \U891/U1117_0_/nd , \U891/U1117_0_/n2 , \U891/U1117_1_/nr , 
        \U891/U1117_1_/nd , \U891/U1117_1_/n2 , \U891/U1117_2_/nr , 
        \U891/U1117_2_/nd , \U891/U1117_2_/n2 , \U891/U1117_3_/nr , 
        \U891/U1117_3_/nd , \U891/U1117_3_/n2 , \U886/nack , \U886/acka , 
        \U886/ackb , \U886/reset , \U886/U1128/nb , \U886/U1128/na , 
        \U886/U1127/n5 , \U886/U1127/n1 , \U886/U1127/n2 , \U886/U1127/n3 , 
        \U886/U1127/n4 , \U886/U1118_0_/nr , \U886/U1118_0_/nd , 
        \U886/U1118_0_/n2 , \U886/U1118_1_/nr , \U886/U1118_1_/nd , 
        \U886/U1118_1_/n2 , \U886/U1118_2_/nr , \U886/U1118_2_/nd , 
        \U886/U1118_2_/n2 , \U886/U1118_3_/nr , \U886/U1118_3_/nd , 
        \U886/U1118_3_/n2 , \U886/U1117_0_/nr , \U886/U1117_0_/nd , 
        \U886/U1117_0_/n2 , \U886/U1117_1_/nr , \U886/U1117_1_/nd , 
        \U886/U1117_1_/n2 , \U886/U1117_2_/nr , \U886/U1117_2_/nd , 
        \U886/U1117_2_/n2 , \U886/U1117_3_/nr , \U886/U1117_3_/nd , 
        \U886/U1117_3_/n2 , \U884/nack , \U884/acka , \U884/ackb , 
        \U884/reset , \U884/U1128/nb , \U884/U1128/na , \U884/U1127/n5 , 
        \U884/U1127/n1 , \U884/U1127/n2 , \U884/U1127/n3 , \U884/U1127/n4 , 
        \U884/U1118_0_/nr , \U884/U1118_0_/nd , \U884/U1118_0_/n2 , 
        \U884/U1118_1_/nr , \U884/U1118_1_/nd , \U884/U1118_1_/n2 , 
        \U884/U1118_2_/nr , \U884/U1118_2_/nd , \U884/U1118_2_/n2 , 
        \U884/U1118_3_/nr , \U884/U1118_3_/nd , \U884/U1118_3_/n2 , 
        \U884/U1117_0_/nr , \U884/U1117_0_/nd , \U884/U1117_0_/n2 , 
        \U884/U1117_1_/nr , \U884/U1117_1_/nd , \U884/U1117_1_/n2 , 
        \U884/U1117_2_/nr , \U884/U1117_2_/nd , \U884/U1117_2_/n2 , 
        \U884/U1117_3_/nr , \U884/U1117_3_/nd , \U884/U1117_3_/n2 , 
        \U888/naack , \U888/r , \U888/s , \U888/nback , \U888/reset , 
        \U887/naack , \U887/r , \U887/s , \U887/nback , \U887/reset , 
        \U885/naack , \U885/r , \U885/s , \U885/nback , \U885/reset , \U877/x , 
        \U877/y , \U877/reset , \U877/U590/U25/U1/clr , \U877/U590/U25/U1/ob , 
        \U877/U589/U25/U1/clr , \U877/U589/U25/U1/ob , \U877/U588/U25/U1/clr , 
        \U877/U588/U25/U1/ob , \U877/U591/U25/U1/clr , \U877/U591/U25/U1/ob , 
        \U876/x , \U876/y , \U876/reset , \U876/U590/U25/U1/clr , 
        \U876/U590/U25/U1/ob , \U876/U589/U25/U1/clr , \U876/U589/U25/U1/ob , 
        \U876/U588/U25/U1/clr , \U876/U588/U25/U1/ob , \U876/U591/U25/U1/clr , 
        \U876/U591/U25/U1/ob , \U2/x , \U2/y , \U2/reset , 
        \U2/U590/U25/U1/clr , \U2/U590/U25/U1/ob , \U2/U589/U25/U1/clr , 
        \U2/U589/U25/U1/ob , \U2/U588/U25/U1/clr , \U2/U588/U25/U1/ob , 
        \U2/U591/U25/U1/clr , \U2/U591/U25/U1/ob , \U1/x , \U1/y , \U1/reset , 
        \U1/U590/U25/U1/clr , \U1/U590/U25/U1/ob , \U1/U589/U25/U1/clr , 
        \U1/U589/U25/U1/ob , \U1/U588/U25/U1/clr , \U1/U588/U25/U1/ob , 
        \U1/U591/U25/U1/clr , \U1/U591/U25/U1/ob , \U881/nack[1] , 
        \U881/nack[0] , n1;
    buf_2 U897 ( .x(nbReset), .a(nReset) );
    and4_1 \U894/U12  ( .x(eop), .a(ncla), .b(csela), .c(asela), .d(i[4]) );
    inv_1 \U891/U1126/U3  ( .x(\U891/reset ), .a(nbReset) );
    inv_1 \U891/U1139/U3  ( .x(\U891/neopack ), .a(eop) );
    nand3_1 \U891/U1131/U9  ( .x(\U891/iay ), .a(\U891/neopack ), .b(
        \U891/naack[0] ), .c(\U891/naack[1] ) );
    nor3_1 \U891/U1128/U27  ( .x(\U891/U1128/nb ), .a(\U891/reset ), .b(\b[3] 
        ), .c(\b[2] ) );
    nor2_1 \U891/U1128/U26  ( .x(\U891/U1128/na ), .a(\b[1] ), .b(\b[0] ) );
    nand2_2 \U891/U1128/U29  ( .x(\U891/ackb ), .a(\U891/U1128/nb ), .b(
        \U891/U1128/na ) );
    nor2_1 \U891/U1133/U5  ( .x(\U891/naack[0] ), .a(\a[3] ), .b(\a[2] ) );
    nor2_1 \U891/U1108/U5  ( .x(\U891/nack ), .a(\U891/acka ), .b(\U891/ackb )
         );
    nor2_1 \U891/U1134/U5  ( .x(\U891/naack[1] ), .a(\a[1] ), .b(\a[0] ) );
    nor2_2 \U891/U914/U6  ( .x(nia), .a(\U891/iay ), .b(\U891/ackb ) );
    nand2_1 \U891/U1130/U5  ( .x(\U891/acka ), .a(\U891/naack[0] ), .b(
        \U891/naack[1] ) );
    ao222_4 \U891/U1121/U1/U1  ( .x(bsela), .a(\U891/nack ), .b(bsel), .c(
        \U891/nack ), .d(bsela), .e(bsel), .f(bsela) );
    ao222_4 \U891/U1120/U1/U1  ( .x(asela), .a(asel), .b(\U891/nack ), .c(asel
        ), .d(asela), .e(\U891/nack ), .f(asela) );
    nor3_1 \U891/U1118_0_/Unr  ( .x(\U891/U1118_0_/nr ), .a(i[0]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_0_/Und  ( .x(\U891/U1118_0_/nd ), .a(i[0]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_0_/U1  ( .x(\U891/U1118_0_/n2 ), .a(\U891/U1118_0_/n2 ), 
        .b(\U891/U1118_0_/nr ), .c(\U891/U1118_0_/nd ) );
    inv_2 \U891/U1118_0_/U3  ( .x(\a[0] ), .a(\U891/U1118_0_/n2 ) );
    nor3_1 \U891/U1118_1_/Unr  ( .x(\U891/U1118_1_/nr ), .a(i[1]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_1_/Und  ( .x(\U891/U1118_1_/nd ), .a(i[1]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_1_/U1  ( .x(\U891/U1118_1_/n2 ), .a(\U891/U1118_1_/n2 ), 
        .b(\U891/U1118_1_/nr ), .c(\U891/U1118_1_/nd ) );
    inv_2 \U891/U1118_1_/U3  ( .x(\a[1] ), .a(\U891/U1118_1_/n2 ) );
    nor3_1 \U891/U1118_2_/Unr  ( .x(\U891/U1118_2_/nr ), .a(i[2]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_2_/Und  ( .x(\U891/U1118_2_/nd ), .a(i[2]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_2_/U1  ( .x(\U891/U1118_2_/n2 ), .a(\U891/U1118_2_/n2 ), 
        .b(\U891/U1118_2_/nr ), .c(\U891/U1118_2_/nd ) );
    inv_2 \U891/U1118_2_/U3  ( .x(\a[2] ), .a(\U891/U1118_2_/n2 ) );
    nor3_1 \U891/U1118_3_/Unr  ( .x(\U891/U1118_3_/nr ), .a(i[3]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_3_/Und  ( .x(\U891/U1118_3_/nd ), .a(i[3]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_3_/U1  ( .x(\U891/U1118_3_/n2 ), .a(\U891/U1118_3_/n2 ), 
        .b(\U891/U1118_3_/nr ), .c(\U891/U1118_3_/nd ) );
    inv_2 \U891/U1118_3_/U3  ( .x(\a[3] ), .a(\U891/U1118_3_/n2 ) );
    nor3_1 \U891/U1117_0_/Unr  ( .x(\U891/U1117_0_/nr ), .a(i[0]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_0_/Und  ( .x(\U891/U1117_0_/nd ), .a(i[0]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_0_/U1  ( .x(\U891/U1117_0_/n2 ), .a(\U891/U1117_0_/n2 ), 
        .b(\U891/U1117_0_/nr ), .c(\U891/U1117_0_/nd ) );
    inv_2 \U891/U1117_0_/U3  ( .x(\b[0] ), .a(\U891/U1117_0_/n2 ) );
    nor3_1 \U891/U1117_1_/Unr  ( .x(\U891/U1117_1_/nr ), .a(i[1]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_1_/Und  ( .x(\U891/U1117_1_/nd ), .a(i[1]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_1_/U1  ( .x(\U891/U1117_1_/n2 ), .a(\U891/U1117_1_/n2 ), 
        .b(\U891/U1117_1_/nr ), .c(\U891/U1117_1_/nd ) );
    inv_2 \U891/U1117_1_/U3  ( .x(\b[1] ), .a(\U891/U1117_1_/n2 ) );
    nor3_1 \U891/U1117_2_/Unr  ( .x(\U891/U1117_2_/nr ), .a(i[2]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_2_/Und  ( .x(\U891/U1117_2_/nd ), .a(i[2]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_2_/U1  ( .x(\U891/U1117_2_/n2 ), .a(\U891/U1117_2_/n2 ), 
        .b(\U891/U1117_2_/nr ), .c(\U891/U1117_2_/nd ) );
    inv_2 \U891/U1117_2_/U3  ( .x(\b[2] ), .a(\U891/U1117_2_/n2 ) );
    nor3_1 \U891/U1117_3_/Unr  ( .x(\U891/U1117_3_/nr ), .a(i[3]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_3_/Und  ( .x(\U891/U1117_3_/nd ), .a(i[3]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_3_/U1  ( .x(\U891/U1117_3_/n2 ), .a(\U891/U1117_3_/n2 ), 
        .b(\U891/U1117_3_/nr ), .c(\U891/U1117_3_/nd ) );
    inv_2 \U891/U1117_3_/U3  ( .x(\b[3] ), .a(\U891/U1117_3_/n2 ) );
    inv_1 \U886/U1126/U3  ( .x(\U886/reset ), .a(nbReset) );
    nor3_1 \U886/U1128/U27  ( .x(\U886/U1128/nb ), .a(\U886/reset ), .b(\f[3] 
        ), .c(\f[2] ) );
    nor2_1 \U886/U1128/U26  ( .x(\U886/U1128/na ), .a(\f[1] ), .b(\f[0] ) );
    nand2_2 \U886/U1128/U29  ( .x(\U886/ackb ), .a(\U886/U1128/nb ), .b(
        \U886/U1128/na ) );
    nor2_1 \U886/U1108/U5  ( .x(\U886/nack ), .a(\U886/acka ), .b(\U886/ackb )
         );
    nor2_2 \U886/U914/U6  ( .x(nba), .a(\U886/acka ), .b(\U886/ackb ) );
    and4_1 \U886/U1127/U25  ( .x(\U886/U1127/n5 ), .a(\U886/U1127/n1 ), .b(
        \U886/U1127/n2 ), .c(\U886/U1127/n3 ), .d(\U886/U1127/n4 ) );
    inv_1 \U886/U1127/U1  ( .x(\U886/U1127/n1 ), .a(\e[3] ) );
    inv_1 \U886/U1127/U2  ( .x(\U886/U1127/n2 ), .a(\e[2] ) );
    inv_1 \U886/U1127/U3  ( .x(\U886/U1127/n3 ), .a(\e[1] ) );
    inv_1 \U886/U1127/U4  ( .x(\U886/U1127/n4 ), .a(\e[0] ) );
    inv_2 \U886/U1127/U5  ( .x(\U886/acka ), .a(\U886/U1127/n5 ) );
    ao222_2 \U886/U1121/U19/U1/U1  ( .x(fsela), .a(\U886/nack ), .b(fsel), .c(
        \U886/nack ), .d(fsela), .e(fsel), .f(fsela) );
    ao222_2 \U886/U1120/U19/U1/U1  ( .x(esela), .a(esel), .b(\U886/nack ), .c(
        esel), .d(esela), .e(\U886/nack ), .f(esela) );
    nor3_1 \U886/U1118_0_/Unr  ( .x(\U886/U1118_0_/nr ), .a(\b[0] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_0_/Und  ( .x(\U886/U1118_0_/nd ), .a(\b[0] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_0_/U1  ( .x(\U886/U1118_0_/n2 ), .a(\U886/U1118_0_/n2 ), 
        .b(\U886/U1118_0_/nr ), .c(\U886/U1118_0_/nd ) );
    inv_2 \U886/U1118_0_/U3  ( .x(\e[0] ), .a(\U886/U1118_0_/n2 ) );
    nor3_1 \U886/U1118_1_/Unr  ( .x(\U886/U1118_1_/nr ), .a(\b[1] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_1_/Und  ( .x(\U886/U1118_1_/nd ), .a(\b[1] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_1_/U1  ( .x(\U886/U1118_1_/n2 ), .a(\U886/U1118_1_/n2 ), 
        .b(\U886/U1118_1_/nr ), .c(\U886/U1118_1_/nd ) );
    inv_2 \U886/U1118_1_/U3  ( .x(\e[1] ), .a(\U886/U1118_1_/n2 ) );
    nor3_1 \U886/U1118_2_/Unr  ( .x(\U886/U1118_2_/nr ), .a(\b[2] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_2_/Und  ( .x(\U886/U1118_2_/nd ), .a(\b[2] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_2_/U1  ( .x(\U886/U1118_2_/n2 ), .a(\U886/U1118_2_/n2 ), 
        .b(\U886/U1118_2_/nr ), .c(\U886/U1118_2_/nd ) );
    inv_2 \U886/U1118_2_/U3  ( .x(\e[2] ), .a(\U886/U1118_2_/n2 ) );
    nor3_1 \U886/U1118_3_/Unr  ( .x(\U886/U1118_3_/nr ), .a(\b[3] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_3_/Und  ( .x(\U886/U1118_3_/nd ), .a(\b[3] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_3_/U1  ( .x(\U886/U1118_3_/n2 ), .a(\U886/U1118_3_/n2 ), 
        .b(\U886/U1118_3_/nr ), .c(\U886/U1118_3_/nd ) );
    inv_2 \U886/U1118_3_/U3  ( .x(\e[3] ), .a(\U886/U1118_3_/n2 ) );
    nor3_1 \U886/U1117_0_/Unr  ( .x(\U886/U1117_0_/nr ), .a(\b[0] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_0_/Und  ( .x(\U886/U1117_0_/nd ), .a(\b[0] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_0_/U1  ( .x(\U886/U1117_0_/n2 ), .a(\U886/U1117_0_/n2 ), 
        .b(\U886/U1117_0_/nr ), .c(\U886/U1117_0_/nd ) );
    inv_2 \U886/U1117_0_/U3  ( .x(\f[0] ), .a(\U886/U1117_0_/n2 ) );
    nor3_1 \U886/U1117_1_/Unr  ( .x(\U886/U1117_1_/nr ), .a(\b[1] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_1_/Und  ( .x(\U886/U1117_1_/nd ), .a(\b[1] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_1_/U1  ( .x(\U886/U1117_1_/n2 ), .a(\U886/U1117_1_/n2 ), 
        .b(\U886/U1117_1_/nr ), .c(\U886/U1117_1_/nd ) );
    inv_2 \U886/U1117_1_/U3  ( .x(\f[1] ), .a(\U886/U1117_1_/n2 ) );
    nor3_1 \U886/U1117_2_/Unr  ( .x(\U886/U1117_2_/nr ), .a(\b[2] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_2_/Und  ( .x(\U886/U1117_2_/nd ), .a(\b[2] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_2_/U1  ( .x(\U886/U1117_2_/n2 ), .a(\U886/U1117_2_/n2 ), 
        .b(\U886/U1117_2_/nr ), .c(\U886/U1117_2_/nd ) );
    inv_2 \U886/U1117_2_/U3  ( .x(\f[2] ), .a(\U886/U1117_2_/n2 ) );
    nor3_1 \U886/U1117_3_/Unr  ( .x(\U886/U1117_3_/nr ), .a(\b[3] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_3_/Und  ( .x(\U886/U1117_3_/nd ), .a(\b[3] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_3_/U1  ( .x(\U886/U1117_3_/n2 ), .a(\U886/U1117_3_/n2 ), 
        .b(\U886/U1117_3_/nr ), .c(\U886/U1117_3_/nd ) );
    inv_2 \U886/U1117_3_/U3  ( .x(\f[3] ), .a(\U886/U1117_3_/n2 ) );
    inv_1 \U884/U1126/U3  ( .x(\U884/reset ), .a(nbReset) );
    nor3_1 \U884/U1128/U27  ( .x(\U884/U1128/nb ), .a(\U884/reset ), .b(\d[3] 
        ), .c(\d[2] ) );
    nor2_1 \U884/U1128/U26  ( .x(\U884/U1128/na ), .a(\d[1] ), .b(\d[0] ) );
    nand2_2 \U884/U1128/U29  ( .x(\U884/ackb ), .a(\U884/U1128/nb ), .b(
        \U884/U1128/na ) );
    nor2_1 \U884/U1108/U5  ( .x(\U884/nack ), .a(\U884/acka ), .b(\U884/ackb )
         );
    nor2_2 \U884/U914/U6  ( .x(naa), .a(\U884/acka ), .b(\U884/ackb ) );
    and4_1 \U884/U1127/U25  ( .x(\U884/U1127/n5 ), .a(\U884/U1127/n1 ), .b(
        \U884/U1127/n2 ), .c(\U884/U1127/n3 ), .d(\U884/U1127/n4 ) );
    inv_1 \U884/U1127/U1  ( .x(\U884/U1127/n1 ), .a(\c[3] ) );
    inv_1 \U884/U1127/U2  ( .x(\U884/U1127/n2 ), .a(\c[2] ) );
    inv_1 \U884/U1127/U3  ( .x(\U884/U1127/n3 ), .a(\c[1] ) );
    inv_1 \U884/U1127/U4  ( .x(\U884/U1127/n4 ), .a(\c[0] ) );
    inv_2 \U884/U1127/U5  ( .x(\U884/acka ), .a(\U884/U1127/n5 ) );
    ao222_2 \U884/U1121/U19/U1/U1  ( .x(dsela), .a(\U884/nack ), .b(dsel), .c(
        \U884/nack ), .d(dsela), .e(dsel), .f(dsela) );
    ao222_2 \U884/U1120/U19/U1/U1  ( .x(csela), .a(csel), .b(\U884/nack ), .c(
        csel), .d(csela), .e(\U884/nack ), .f(csela) );
    nor3_1 \U884/U1118_0_/Unr  ( .x(\U884/U1118_0_/nr ), .a(\a[0] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_0_/Und  ( .x(\U884/U1118_0_/nd ), .a(\a[0] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_0_/U1  ( .x(\U884/U1118_0_/n2 ), .a(\U884/U1118_0_/n2 ), 
        .b(\U884/U1118_0_/nr ), .c(\U884/U1118_0_/nd ) );
    inv_2 \U884/U1118_0_/U3  ( .x(\c[0] ), .a(\U884/U1118_0_/n2 ) );
    nor3_1 \U884/U1118_1_/Unr  ( .x(\U884/U1118_1_/nr ), .a(\a[1] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_1_/Und  ( .x(\U884/U1118_1_/nd ), .a(\a[1] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_1_/U1  ( .x(\U884/U1118_1_/n2 ), .a(\U884/U1118_1_/n2 ), 
        .b(\U884/U1118_1_/nr ), .c(\U884/U1118_1_/nd ) );
    inv_2 \U884/U1118_1_/U3  ( .x(\c[1] ), .a(\U884/U1118_1_/n2 ) );
    nor3_1 \U884/U1118_2_/Unr  ( .x(\U884/U1118_2_/nr ), .a(\a[2] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_2_/Und  ( .x(\U884/U1118_2_/nd ), .a(\a[2] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_2_/U1  ( .x(\U884/U1118_2_/n2 ), .a(\U884/U1118_2_/n2 ), 
        .b(\U884/U1118_2_/nr ), .c(\U884/U1118_2_/nd ) );
    inv_2 \U884/U1118_2_/U3  ( .x(\c[2] ), .a(\U884/U1118_2_/n2 ) );
    nor3_1 \U884/U1118_3_/Unr  ( .x(\U884/U1118_3_/nr ), .a(\a[3] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_3_/Und  ( .x(\U884/U1118_3_/nd ), .a(\a[3] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_3_/U1  ( .x(\U884/U1118_3_/n2 ), .a(\U884/U1118_3_/n2 ), 
        .b(\U884/U1118_3_/nr ), .c(\U884/U1118_3_/nd ) );
    inv_2 \U884/U1118_3_/U3  ( .x(\c[3] ), .a(\U884/U1118_3_/n2 ) );
    nor3_1 \U884/U1117_0_/Unr  ( .x(\U884/U1117_0_/nr ), .a(\a[0] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_0_/Und  ( .x(\U884/U1117_0_/nd ), .a(\a[0] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_0_/U1  ( .x(\U884/U1117_0_/n2 ), .a(\U884/U1117_0_/n2 ), 
        .b(\U884/U1117_0_/nr ), .c(\U884/U1117_0_/nd ) );
    inv_2 \U884/U1117_0_/U3  ( .x(\d[0] ), .a(\U884/U1117_0_/n2 ) );
    nor3_1 \U884/U1117_1_/Unr  ( .x(\U884/U1117_1_/nr ), .a(\a[1] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_1_/Und  ( .x(\U884/U1117_1_/nd ), .a(\a[1] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_1_/U1  ( .x(\U884/U1117_1_/n2 ), .a(\U884/U1117_1_/n2 ), 
        .b(\U884/U1117_1_/nr ), .c(\U884/U1117_1_/nd ) );
    inv_2 \U884/U1117_1_/U3  ( .x(\d[1] ), .a(\U884/U1117_1_/n2 ) );
    nor3_1 \U884/U1117_2_/Unr  ( .x(\U884/U1117_2_/nr ), .a(\a[2] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_2_/Und  ( .x(\U884/U1117_2_/nd ), .a(\a[2] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_2_/U1  ( .x(\U884/U1117_2_/n2 ), .a(\U884/U1117_2_/n2 ), 
        .b(\U884/U1117_2_/nr ), .c(\U884/U1117_2_/nd ) );
    inv_2 \U884/U1117_2_/U3  ( .x(\d[2] ), .a(\U884/U1117_2_/n2 ) );
    nor3_1 \U884/U1117_3_/Unr  ( .x(\U884/U1117_3_/nr ), .a(\a[3] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_3_/Und  ( .x(\U884/U1117_3_/nd ), .a(\a[3] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_3_/U1  ( .x(\U884/U1117_3_/n2 ), .a(\U884/U1117_3_/n2 ), 
        .b(\U884/U1117_3_/nr ), .c(\U884/U1117_3_/nd ) );
    inv_2 \U884/U1117_3_/U3  ( .x(\d[3] ), .a(\U884/U1117_3_/n2 ) );
    nand2_1 \U888/U1128/U5  ( .x(\U888/s ), .a(\U888/r ), .b(\U888/nback ) );
    nand2_1 \U888/U1103/U5  ( .x(\U888/r ), .a(\U888/naack ), .b(\U888/s ) );
    inv_1 \U888/U1111/U3  ( .x(\U888/reset ), .a(nbReset) );
    inv_1 \U888/U1112/U3  ( .x(\U888/naack ), .a(esela) );
    nor2_1 \U888/U1127/U5  ( .x(\U888/nback ), .a(fsela), .b(\U888/reset ) );
    and2_2 \U888/U1129/U8  ( .x(esel), .a(\U888/nback ), .b(\U888/s ) );
    and2_2 \U888/U1124/U8  ( .x(fsel), .a(\U888/r ), .b(\U888/naack ) );
    nand2_1 \U887/U1128/U5  ( .x(\U887/s ), .a(\U887/r ), .b(\U887/nback ) );
    nand2_1 \U887/U1103/U5  ( .x(\U887/r ), .a(\U887/naack ), .b(\U887/s ) );
    inv_1 \U887/U1111/U3  ( .x(\U887/reset ), .a(nbReset) );
    inv_1 \U887/U1112/U3  ( .x(\U887/naack ), .a(csela) );
    nor2_1 \U887/U1127/U5  ( .x(\U887/nback ), .a(dsela), .b(\U887/reset ) );
    and2_2 \U887/U1129/U8  ( .x(csel), .a(\U887/nback ), .b(\U887/s ) );
    and2_2 \U887/U1124/U8  ( .x(dsel), .a(\U887/r ), .b(\U887/naack ) );
    nand2_1 \U885/U1128/U5  ( .x(\U885/s ), .a(\U885/r ), .b(\U885/nback ) );
    nand2_1 \U885/U1103/U5  ( .x(\U885/r ), .a(\U885/naack ), .b(\U885/s ) );
    inv_1 \U885/U1111/U3  ( .x(\U885/reset ), .a(nbReset) );
    inv_1 \U885/U1112/U3  ( .x(\U885/naack ), .a(asela) );
    nor2_1 \U885/U1127/U5  ( .x(\U885/nback ), .a(bsela), .b(\U885/reset ) );
    and2_2 \U885/U1129/U8  ( .x(asel), .a(\U885/nback ), .b(\U885/s ) );
    and2_2 \U885/U1124/U8  ( .x(bsel), .a(\U885/r ), .b(\U885/naack ) );
    nor3_1 \U877/U594/U7  ( .x(\U877/x ), .a(ol[7]), .b(\U877/reset ), .c(oh
        [7]) );
    nor3_1 \U877/U593/U7  ( .x(\U877/y ), .a(ol[6]), .b(\U877/reset ), .c(oh
        [6]) );
    inv_1 \U877/U604/U3  ( .x(\U877/reset ), .a(nbReset) );
    oa31_1 \U877/U590/U25/U1/Uclr  ( .x(\U877/U590/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[1] ), .d(oh[6]) );
    oaoi211_1 \U877/U590/U25/U1/Uaoi  ( .x(\U877/U590/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[1] ), .c(n1), .d(\U877/U590/U25/U1/clr ) );
    inv_2 \U877/U590/U25/U1/Ui  ( .x(oh[6]), .a(\U877/U590/U25/U1/ob ) );
    oa31_1 \U877/U589/U25/U1/Uclr  ( .x(\U877/U589/U25/U1/clr ), .a(net135), 
        .b(\cl[1] ), .c(\cl[0] ), .d(ol[7]) );
    oaoi211_1 \U877/U589/U25/U1/Uaoi  ( .x(\U877/U589/U25/U1/ob ), .a(\cl[1] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U589/U25/U1/clr ) );
    inv_2 \U877/U589/U25/U1/Ui  ( .x(ol[7]), .a(\U877/U589/U25/U1/ob ) );
    oa31_1 \U877/U588/U25/U1/Uclr  ( .x(\U877/U588/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[2] ), .d(oh[7]) );
    oaoi211_1 \U877/U588/U25/U1/Uaoi  ( .x(\U877/U588/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[2] ), .c(n1), .d(\U877/U588/U25/U1/clr ) );
    inv_2 \U877/U588/U25/U1/Ui  ( .x(oh[7]), .a(\U877/U588/U25/U1/ob ) );
    oa31_1 \U877/U591/U25/U1/Uclr  ( .x(\U877/U591/U25/U1/clr ), .a(net135), 
        .b(\cl[2] ), .c(\cl[0] ), .d(ol[6]) );
    oaoi211_1 \U877/U591/U25/U1/Uaoi  ( .x(\U877/U591/U25/U1/ob ), .a(\cl[2] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U591/U25/U1/clr ) );
    inv_2 \U877/U591/U25/U1/Ui  ( .x(ol[6]), .a(\U877/U591/U25/U1/ob ) );
    ao222_2 \U877/U592/U19/U1/U1  ( .x(ncla), .a(\U877/x ), .b(\U877/y ), .c(
        \U877/x ), .d(ncla), .e(\U877/y ), .f(ncla) );
    nor3_1 \U876/U594/U7  ( .x(\U876/x ), .a(ol[3]), .b(\U876/reset ), .c(oh
        [3]) );
    nor3_1 \U876/U593/U7  ( .x(\U876/y ), .a(ol[2]), .b(\U876/reset ), .c(oh
        [2]) );
    inv_1 \U876/U604/U3  ( .x(\U876/reset ), .a(nbReset) );
    oa31_1 \U876/U590/U25/U1/Uclr  ( .x(\U876/U590/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[1] ), .d(oh[2]) );
    oaoi211_1 \U876/U590/U25/U1/Uaoi  ( .x(\U876/U590/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[1] ), .c(n1), .d(\U876/U590/U25/U1/clr ) );
    inv_2 \U876/U590/U25/U1/Ui  ( .x(oh[2]), .a(\U876/U590/U25/U1/ob ) );
    oa31_1 \U876/U589/U25/U1/Uclr  ( .x(\U876/U589/U25/U1/clr ), .a(net135), 
        .b(\d[1] ), .c(\d[0] ), .d(ol[3]) );
    oaoi211_1 \U876/U589/U25/U1/Uaoi  ( .x(\U876/U589/U25/U1/ob ), .a(\d[1] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U589/U25/U1/clr ) );
    inv_2 \U876/U589/U25/U1/Ui  ( .x(ol[3]), .a(\U876/U589/U25/U1/ob ) );
    oa31_1 \U876/U588/U25/U1/Uclr  ( .x(\U876/U588/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[2] ), .d(oh[3]) );
    oaoi211_1 \U876/U588/U25/U1/Uaoi  ( .x(\U876/U588/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[2] ), .c(n1), .d(\U876/U588/U25/U1/clr ) );
    inv_2 \U876/U588/U25/U1/Ui  ( .x(oh[3]), .a(\U876/U588/U25/U1/ob ) );
    oa31_1 \U876/U591/U25/U1/Uclr  ( .x(\U876/U591/U25/U1/clr ), .a(net135), 
        .b(\d[2] ), .c(\d[0] ), .d(ol[2]) );
    oaoi211_1 \U876/U591/U25/U1/Uaoi  ( .x(\U876/U591/U25/U1/ob ), .a(\d[2] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U591/U25/U1/clr ) );
    inv_2 \U876/U591/U25/U1/Ui  ( .x(ol[2]), .a(\U876/U591/U25/U1/ob ) );
    ao222_2 \U876/U592/U19/U1/U1  ( .x(nda), .a(\U876/x ), .b(\U876/y ), .c(
        \U876/x ), .d(nda), .e(\U876/y ), .f(nda) );
    nor3_1 \U2/U594/U7  ( .x(\U2/x ), .a(ol[1]), .b(\U2/reset ), .c(oh[1]) );
    nor3_1 \U2/U593/U7  ( .x(\U2/y ), .a(ol[0]), .b(\U2/reset ), .c(oh[0]) );
    inv_1 \U2/U604/U3  ( .x(\U2/reset ), .a(nbReset) );
    oa31_1 \U2/U590/U25/U1/Uclr  ( .x(\U2/U590/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[1] ), .d(oh[0]) );
    oaoi211_1 \U2/U590/U25/U1/Uaoi  ( .x(\U2/U590/U25/U1/ob ), .a(\f[3] ), .b(
        \f[1] ), .c(n1), .d(\U2/U590/U25/U1/clr ) );
    inv_2 \U2/U590/U25/U1/Ui  ( .x(oh[0]), .a(\U2/U590/U25/U1/ob ) );
    oa31_1 \U2/U589/U25/U1/Uclr  ( .x(\U2/U589/U25/U1/clr ), .a(net135), .b(
        \f[1] ), .c(\f[0] ), .d(ol[1]) );
    oaoi211_1 \U2/U589/U25/U1/Uaoi  ( .x(\U2/U589/U25/U1/ob ), .a(\f[1] ), .b(
        \f[0] ), .c(n1), .d(\U2/U589/U25/U1/clr ) );
    inv_2 \U2/U589/U25/U1/Ui  ( .x(ol[1]), .a(\U2/U589/U25/U1/ob ) );
    oa31_1 \U2/U588/U25/U1/Uclr  ( .x(\U2/U588/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[2] ), .d(oh[1]) );
    oaoi211_1 \U2/U588/U25/U1/Uaoi  ( .x(\U2/U588/U25/U1/ob ), .a(\f[3] ), .b(
        \f[2] ), .c(n1), .d(\U2/U588/U25/U1/clr ) );
    inv_2 \U2/U588/U25/U1/Ui  ( .x(oh[1]), .a(\U2/U588/U25/U1/ob ) );
    oa31_1 \U2/U591/U25/U1/Uclr  ( .x(\U2/U591/U25/U1/clr ), .a(net135), .b(
        \f[2] ), .c(\f[0] ), .d(ol[0]) );
    oaoi211_1 \U2/U591/U25/U1/Uaoi  ( .x(\U2/U591/U25/U1/ob ), .a(\f[2] ), .b(
        \f[0] ), .c(n1), .d(\U2/U591/U25/U1/clr ) );
    inv_2 \U2/U591/U25/U1/Ui  ( .x(ol[0]), .a(\U2/U591/U25/U1/ob ) );
    ao222_2 \U2/U592/U19/U1/U1  ( .x(nfa), .a(\U2/x ), .b(\U2/y ), .c(\U2/x ), 
        .d(nfa), .e(\U2/y ), .f(nfa) );
    nor3_1 \U1/U594/U7  ( .x(\U1/x ), .a(ol[5]), .b(\U1/reset ), .c(oh[5]) );
    nor3_1 \U1/U593/U7  ( .x(\U1/y ), .a(ol[4]), .b(\U1/reset ), .c(oh[4]) );
    inv_1 \U1/U604/U3  ( .x(\U1/reset ), .a(nbReset) );
    oa31_1 \U1/U590/U25/U1/Uclr  ( .x(\U1/U590/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[1] ), .d(oh[4]) );
    oaoi211_1 \U1/U590/U25/U1/Uaoi  ( .x(\U1/U590/U25/U1/ob ), .a(\e[3] ), .b(
        \e[1] ), .c(n1), .d(\U1/U590/U25/U1/clr ) );
    inv_2 \U1/U590/U25/U1/Ui  ( .x(oh[4]), .a(\U1/U590/U25/U1/ob ) );
    oa31_1 \U1/U589/U25/U1/Uclr  ( .x(\U1/U589/U25/U1/clr ), .a(net135), .b(
        \e[1] ), .c(\e[0] ), .d(ol[5]) );
    oaoi211_1 \U1/U589/U25/U1/Uaoi  ( .x(\U1/U589/U25/U1/ob ), .a(\e[1] ), .b(
        \e[0] ), .c(n1), .d(\U1/U589/U25/U1/clr ) );
    inv_2 \U1/U589/U25/U1/Ui  ( .x(ol[5]), .a(\U1/U589/U25/U1/ob ) );
    oa31_1 \U1/U588/U25/U1/Uclr  ( .x(\U1/U588/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[2] ), .d(oh[5]) );
    oaoi211_1 \U1/U588/U25/U1/Uaoi  ( .x(\U1/U588/U25/U1/ob ), .a(\e[3] ), .b(
        \e[2] ), .c(n1), .d(\U1/U588/U25/U1/clr ) );
    inv_2 \U1/U588/U25/U1/Ui  ( .x(oh[5]), .a(\U1/U588/U25/U1/ob ) );
    oa31_1 \U1/U591/U25/U1/Uclr  ( .x(\U1/U591/U25/U1/clr ), .a(net135), .b(
        \e[2] ), .c(\e[0] ), .d(ol[4]) );
    oaoi211_1 \U1/U591/U25/U1/Uaoi  ( .x(\U1/U591/U25/U1/ob ), .a(\e[2] ), .b(
        \e[0] ), .c(n1), .d(\U1/U591/U25/U1/clr ) );
    inv_2 \U1/U591/U25/U1/Ui  ( .x(ol[4]), .a(\U1/U591/U25/U1/ob ) );
    ao222_2 \U1/U592/U19/U1/U1  ( .x(nea), .a(\U1/x ), .b(\U1/y ), .c(\U1/x ), 
        .d(nea), .e(\U1/y ), .f(nea) );
    and3_4 \U881/U20/U9  ( .x(nca), .a(\U881/nack[1] ), .b(\U881/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U881/U18/U5  ( .x(\U881/nack[0] ), .a(\cl[3] ), .b(\cl[0] ) );
    nor2_1 \U881/U19/U5  ( .x(\U881/nack[1] ), .a(\cl[1] ), .b(\cl[2] ) );
    ao222_2 \U881/U15_0_/U19/U1/U1  ( .x(\cl[0] ), .a(\c[0] ), .b(ncla), .c(
        \c[0] ), .d(\cl[0] ), .e(ncla), .f(\cl[0] ) );
    ao222_2 \U881/U15_1_/U19/U1/U1  ( .x(\cl[1] ), .a(\c[1] ), .b(ncla), .c(
        \c[1] ), .d(\cl[1] ), .e(ncla), .f(\cl[1] ) );
    ao222_2 \U881/U15_2_/U19/U1/U1  ( .x(\cl[2] ), .a(\c[2] ), .b(ncla), .c(
        \c[2] ), .d(\cl[2] ), .e(ncla), .f(\cl[2] ) );
    ao222_2 \U881/U15_3_/U19/U1/U1  ( .x(\cl[3] ), .a(\c[3] ), .b(ncla), .c(
        \c[3] ), .d(\cl[3] ), .e(ncla), .f(\cl[3] ) );
    and2_5 U1 ( .x(n1), .a(nbReset), .b(noa) );
    and2_3 U2 ( .x(net135), .a(nbReset), .b(noa) );
endmodule


module chain_dr2fr_byte_5 ( eop_ack, ia, o, eop, ih, il, nReset, noa );
output [4:0] o;
input  [7:0] ih;
input  [7:0] il;
input  eop, nReset, noa;
output eop_ack, ia;
    wire eop_pass, nhighack, nlowack, \twobitack[2] , \twobitack[3] , 
        \twobitack[0] , \twobitack[1] , xsel, ysel, nxa, nyla, nbReset, nya, 
        \y[3] , \y[2] , \y[1] , \y[0] , \yl[3] , \yl[2] , \yl[1] , \yl[0] , 
        \cdh[0] , \cdh[1] , \cdl[0] , \cdl[1] , net193, \cdh[2] , \cdh[3] , 
        \cdl[2] , \cdl[3] , net195, bsel, dsel, nba, bg, nda, dg, asel, csel, 
        naa, ag, nca, cg, \d[3] , \d[2] , \d[1] , \d[0] , \b[3] , \b[2] , 
        \b[1] , \b[0] , \x[3] , \x[2] , \x[1] , \x[0] , \c[3] , \c[2] , \c[1] , 
        \c[0] , \a[3] , \a[2] , \a[1] , \a[0] , net194, net199, \U1018/Z , 
        \U1270/net190 , \U1270/net191 , \U1270/net192 , \U1270/net189 , 
        \U1270/U1141/Z , \U1268/net190 , \U1268/net191 , \U1268/net192 , 
        \U1268/net189 , \U1268/U1141/Z , \U1224/nack[0] , \U1224/nack[1] , 
        \U1224/net4 , \U1224/U1125/U28/U1/clr , \U1224/U1125/U28/U1/set , 
        \U1224/U1122/U28/U1/clr , \U1224/U1122/U28/U1/set , 
        \U1224/U916_0_/U25/U1/clr , \U1224/U916_0_/U25/U1/ob , 
        \U1224/U916_1_/U25/U1/clr , \U1224/U916_1_/U25/U1/ob , 
        \U1224/U916_2_/U25/U1/clr , \U1224/U916_2_/U25/U1/ob , 
        \U1224/U916_3_/U25/U1/clr , \U1224/U916_3_/U25/U1/ob , \U1209/nack[0] , 
        \U1209/nack[1] , \U1209/net4 , \U1209/U1125/U28/U1/clr , 
        \U1209/U1125/U28/U1/set , \U1209/U1122/U28/U1/clr , 
        \U1209/U1122/U28/U1/set , \U1209/U916_0_/U25/U1/clr , 
        \U1209/U916_0_/U25/U1/ob , \U1209/U916_1_/U25/U1/clr , 
        \U1209/U916_1_/U25/U1/ob , \U1209/U916_2_/U25/U1/clr , 
        \U1209/U916_2_/U25/U1/ob , \U1209/U916_3_/U25/U1/clr , 
        \U1209/U916_3_/U25/U1/ob , \U1213/nack[0] , \U1213/nack[1] , 
        \U1213/net4 , \U1213/U1125/U28/U1/clr , \U1213/U1125/U28/U1/set , 
        \U1213/U1122/U28/U1/clr , \U1213/U1122/U28/U1/set , 
        \U1213/U916_0_/U25/U1/clr , \U1213/U916_0_/U25/U1/ob , 
        \U1213/U916_1_/U25/U1/clr , \U1213/U916_1_/U25/U1/ob , 
        \U1213/U916_2_/U25/U1/clr , \U1213/U916_2_/U25/U1/ob , 
        \U1213/U916_3_/U25/U1/clr , \U1213/U916_3_/U25/U1/ob , \U1296/ng , 
        \U1296/U1384/Z , \U1296/U1386/U25/U1/clr , \U1296/U1386/U25/U1/ob , 
        \U1298/ng , \U1298/U1384/Z , \U1298/U1386/U25/U1/clr , 
        \U1298/U1386/U25/U1/ob , \U1306/ng , \U1306/U1384/Z , 
        \U1306/U1386/U25/U1/clr , \U1306/U1386/U25/U1/ob , \U1295/ng , 
        \U1295/U1384/Z , \U1295/U1386/U25/U1/clr , \U1295/U1386/U25/U1/ob , 
        \U1297/s , \U1297/nback , \U1297/r , \U1297/naack , \U1297/reset , 
        \U1297/U1128/U28/U1/clr , \U1297/U1128/U28/U1/set , 
        \U1297/U1127/U28/U1/clr , \U1297/U1127/U28/U1/set , \U1300/s , 
        \U1300/nback , \U1300/r , \U1300/naack , \U1300/reset , 
        \U1300/U1128/U28/U1/clr , \U1300/U1128/U28/U1/set , 
        \U1300/U1127/U28/U1/clr , \U1300/U1127/U28/U1/set , \U1289/bnreset , 
        \U1289/U1150/U28/U1/clr , \U1289/U1150/U28/U1/set , 
        \U1289/U1152/U28/U1/clr , \U1289/U1152/U28/U1/set , 
        \U1289/U1149/U28/U1/clr , \U1289/U1149/U28/U1/set , 
        \U1289/U1151/U28/U1/clr , \U1289/U1151/U28/U1/set , 
        \U1289/U1148/net190 , \U1289/U1148/net191 , \U1289/U1148/net192 , 
        \U1289/U1148/net189 , \U1289/U1148/U1141/Z , \U1271/bnreset , 
        \U1271/U1150/U28/U1/clr , \U1271/U1150/U28/U1/set , 
        \U1271/U1152/U28/U1/clr , \U1271/U1152/U28/U1/set , 
        \U1271/U1149/U28/U1/clr , \U1271/U1149/U28/U1/set , 
        \U1271/U1151/U28/U1/clr , \U1271/U1151/U28/U1/set , 
        \U1271/U1148/net190 , \U1271/U1148/net191 , \U1271/U1148/net192 , 
        \U1271/U1148/net189 , \U1271/U1148/U1141/Z , \U1225/naack , \U1225/r , 
        \U1225/s , \U1225/nback , \U1225/reset , \U1308/nack[1] , 
        \U1308/nack[0] ;
    assign o[4] = eop_ack;
    buf_2 U1231 ( .x(nbReset), .a(nReset) );
    and3_1 \U1194/U9  ( .x(eop_pass), .a(nxa), .b(naa), .c(eop) );
    ao222_1 \U1301/U18/U1/U1  ( .x(nlowack), .a(\twobitack[0] ), .b(
        \twobitack[1] ), .c(\twobitack[0] ), .d(nlowack), .e(\twobitack[1] ), 
        .f(nlowack) );
    ao222_1 \U1302/U18/U1/U1  ( .x(nhighack), .a(\twobitack[2] ), .b(
        \twobitack[3] ), .c(\twobitack[2] ), .d(nhighack), .e(\twobitack[3] ), 
        .f(nhighack) );
    aoi222_1 \U1018/U30/U1  ( .x(ia), .a(nhighack), .b(nlowack), .c(nhighack), 
        .d(\U1018/Z ), .e(nlowack), .f(\U1018/Z ) );
    inv_1 \U1018/U30/Uinv  ( .x(\U1018/Z ), .a(ia) );
    ao222_2 \U1038/U19/U1/U1  ( .x(eop_ack), .a(eop_pass), .b(noa), .c(
        eop_pass), .d(eop_ack), .e(noa), .f(eop_ack) );
    inv_1 \U1270/U1147/U3  ( .x(\U1270/net189 ), .a(nbReset) );
    nor2_1 \U1270/U582/U5  ( .x(\U1270/net192 ), .a(il[4]), .b(ih[4]) );
    nor2_1 \U1270/U580/U5  ( .x(\U1270/net191 ), .a(il[5]), .b(ih[5]) );
    nor2_2 \U1270/U1146/U6  ( .x(net199), .a(\U1270/net190 ), .b(
        \U1270/net189 ) );
    aoi222_1 \U1270/U1141/U30/U1  ( .x(\U1270/net190 ), .a(\U1270/net191 ), 
        .b(\U1270/net192 ), .c(\U1270/net191 ), .d(\U1270/U1141/Z ), .e(
        \U1270/net192 ), .f(\U1270/U1141/Z ) );
    inv_1 \U1270/U1141/U30/Uinv  ( .x(\U1270/U1141/Z ), .a(\U1270/net190 ) );
    inv_1 \U1268/U1147/U3  ( .x(\U1268/net189 ), .a(nbReset) );
    nor2_1 \U1268/U582/U5  ( .x(\U1268/net192 ), .a(il[6]), .b(ih[6]) );
    nor2_1 \U1268/U580/U5  ( .x(\U1268/net191 ), .a(il[7]), .b(ih[7]) );
    nor2_2 \U1268/U1146/U6  ( .x(net194), .a(\U1268/net190 ), .b(
        \U1268/net189 ) );
    aoi222_1 \U1268/U1141/U30/U1  ( .x(\U1268/net190 ), .a(\U1268/net191 ), 
        .b(\U1268/net192 ), .c(\U1268/net191 ), .d(\U1268/U1141/Z ), .e(
        \U1268/net192 ), .f(\U1268/U1141/Z ) );
    inv_1 \U1268/U1141/U30/Uinv  ( .x(\U1268/U1141/Z ), .a(\U1268/net190 ) );
    nor2_1 \U1224/U1128/U5  ( .x(\U1224/nack[0] ), .a(\x[3] ), .b(\x[2] ) );
    nor3_1 \U1224/U1127/U7  ( .x(\U1224/nack[1] ), .a(\x[1] ), .b(\U1224/net4 
        ), .c(\x[0] ) );
    inv_1 \U1224/U907/U3  ( .x(\U1224/net4 ), .a(nbReset) );
    aoai211_1 \U1224/U1125/U28/U1/U1  ( .x(\U1224/U1125/U28/U1/clr ), .a(
        \U1224/nack[1] ), .b(\U1224/nack[0] ), .c(asel), .d(naa) );
    nand3_1 \U1224/U1125/U28/U1/U2  ( .x(\U1224/U1125/U28/U1/set ), .a(asel), 
        .b(\U1224/nack[1] ), .c(\U1224/nack[0] ) );
    nand2_2 \U1224/U1125/U28/U1/U3  ( .x(naa), .a(\U1224/U1125/U28/U1/clr ), 
        .b(\U1224/U1125/U28/U1/set ) );
    aoai211_1 \U1224/U1122/U28/U1/U1  ( .x(\U1224/U1122/U28/U1/clr ), .a(
        \U1224/nack[0] ), .b(\U1224/nack[1] ), .c(csel), .d(nca) );
    nand3_1 \U1224/U1122/U28/U1/U2  ( .x(\U1224/U1122/U28/U1/set ), .a(csel), 
        .b(\U1224/nack[0] ), .c(\U1224/nack[1] ) );
    nand2_2 \U1224/U1122/U28/U1/U3  ( .x(nca), .a(\U1224/U1122/U28/U1/clr ), 
        .b(\U1224/U1122/U28/U1/set ) );
    oa31_1 \U1224/U916_0_/U25/U1/Uclr  ( .x(\U1224/U916_0_/U25/U1/clr ), .a(
        nxa), .b(\a[0] ), .c(\c[0] ), .d(\x[0] ) );
    oaoi211_1 \U1224/U916_0_/U25/U1/Uaoi  ( .x(\U1224/U916_0_/U25/U1/ob ), .a(
        \a[0] ), .b(\c[0] ), .c(nxa), .d(\U1224/U916_0_/U25/U1/clr ) );
    inv_2 \U1224/U916_0_/U25/U1/Ui  ( .x(\x[0] ), .a(\U1224/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_1_/U25/U1/Uclr  ( .x(\U1224/U916_1_/U25/U1/clr ), .a(
        nxa), .b(\a[1] ), .c(\c[1] ), .d(\x[1] ) );
    oaoi211_1 \U1224/U916_1_/U25/U1/Uaoi  ( .x(\U1224/U916_1_/U25/U1/ob ), .a(
        \a[1] ), .b(\c[1] ), .c(nxa), .d(\U1224/U916_1_/U25/U1/clr ) );
    inv_2 \U1224/U916_1_/U25/U1/Ui  ( .x(\x[1] ), .a(\U1224/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_2_/U25/U1/Uclr  ( .x(\U1224/U916_2_/U25/U1/clr ), .a(
        nxa), .b(\a[2] ), .c(\c[2] ), .d(\x[2] ) );
    oaoi211_1 \U1224/U916_2_/U25/U1/Uaoi  ( .x(\U1224/U916_2_/U25/U1/ob ), .a(
        \a[2] ), .b(\c[2] ), .c(nxa), .d(\U1224/U916_2_/U25/U1/clr ) );
    inv_2 \U1224/U916_2_/U25/U1/Ui  ( .x(\x[2] ), .a(\U1224/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_3_/U25/U1/Uclr  ( .x(\U1224/U916_3_/U25/U1/clr ), .a(
        nxa), .b(\a[3] ), .c(\c[3] ), .d(\x[3] ) );
    oaoi211_1 \U1224/U916_3_/U25/U1/Uaoi  ( .x(\U1224/U916_3_/U25/U1/ob ), .a(
        \a[3] ), .b(\c[3] ), .c(nxa), .d(\U1224/U916_3_/U25/U1/clr ) );
    inv_2 \U1224/U916_3_/U25/U1/Ui  ( .x(\x[3] ), .a(\U1224/U916_3_/U25/U1/ob 
        ) );
    nor2_1 \U1209/U1128/U5  ( .x(\U1209/nack[0] ), .a(o[3]), .b(o[2]) );
    nor3_1 \U1209/U1127/U7  ( .x(\U1209/nack[1] ), .a(o[1]), .b(\U1209/net4 ), 
        .c(o[0]) );
    inv_1 \U1209/U907/U3  ( .x(\U1209/net4 ), .a(nbReset) );
    aoai211_1 \U1209/U1125/U28/U1/U1  ( .x(\U1209/U1125/U28/U1/clr ), .a(
        \U1209/nack[1] ), .b(\U1209/nack[0] ), .c(xsel), .d(nxa) );
    nand3_1 \U1209/U1125/U28/U1/U2  ( .x(\U1209/U1125/U28/U1/set ), .a(xsel), 
        .b(\U1209/nack[1] ), .c(\U1209/nack[0] ) );
    nand2_2 \U1209/U1125/U28/U1/U3  ( .x(nxa), .a(\U1209/U1125/U28/U1/clr ), 
        .b(\U1209/U1125/U28/U1/set ) );
    aoai211_1 \U1209/U1122/U28/U1/U1  ( .x(\U1209/U1122/U28/U1/clr ), .a(
        \U1209/nack[0] ), .b(\U1209/nack[1] ), .c(ysel), .d(nyla) );
    nand3_1 \U1209/U1122/U28/U1/U2  ( .x(\U1209/U1122/U28/U1/set ), .a(ysel), 
        .b(\U1209/nack[0] ), .c(\U1209/nack[1] ) );
    nand2_2 \U1209/U1122/U28/U1/U3  ( .x(nyla), .a(\U1209/U1122/U28/U1/clr ), 
        .b(\U1209/U1122/U28/U1/set ) );
    oa31_1 \U1209/U916_0_/U25/U1/Uclr  ( .x(\U1209/U916_0_/U25/U1/clr ), .a(
        noa), .b(\x[0] ), .c(\yl[0] ), .d(o[0]) );
    oaoi211_1 \U1209/U916_0_/U25/U1/Uaoi  ( .x(\U1209/U916_0_/U25/U1/ob ), .a(
        \x[0] ), .b(\yl[0] ), .c(noa), .d(\U1209/U916_0_/U25/U1/clr ) );
    inv_2 \U1209/U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U1209/U916_0_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_1_/U25/U1/Uclr  ( .x(\U1209/U916_1_/U25/U1/clr ), .a(
        noa), .b(\x[1] ), .c(\yl[1] ), .d(o[1]) );
    oaoi211_1 \U1209/U916_1_/U25/U1/Uaoi  ( .x(\U1209/U916_1_/U25/U1/ob ), .a(
        \x[1] ), .b(\yl[1] ), .c(noa), .d(\U1209/U916_1_/U25/U1/clr ) );
    inv_2 \U1209/U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U1209/U916_1_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_2_/U25/U1/Uclr  ( .x(\U1209/U916_2_/U25/U1/clr ), .a(
        noa), .b(\x[2] ), .c(\yl[2] ), .d(o[2]) );
    oaoi211_1 \U1209/U916_2_/U25/U1/Uaoi  ( .x(\U1209/U916_2_/U25/U1/ob ), .a(
        \x[2] ), .b(\yl[2] ), .c(noa), .d(\U1209/U916_2_/U25/U1/clr ) );
    inv_2 \U1209/U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U1209/U916_2_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_3_/U25/U1/Uclr  ( .x(\U1209/U916_3_/U25/U1/clr ), .a(
        noa), .b(\x[3] ), .c(\yl[3] ), .d(o[3]) );
    oaoi211_1 \U1209/U916_3_/U25/U1/Uaoi  ( .x(\U1209/U916_3_/U25/U1/ob ), .a(
        \x[3] ), .b(\yl[3] ), .c(noa), .d(\U1209/U916_3_/U25/U1/clr ) );
    inv_2 \U1209/U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U1209/U916_3_/U25/U1/ob )
         );
    nor2_1 \U1213/U1128/U5  ( .x(\U1213/nack[0] ), .a(\y[3] ), .b(\y[2] ) );
    nor3_1 \U1213/U1127/U7  ( .x(\U1213/nack[1] ), .a(\y[1] ), .b(\U1213/net4 
        ), .c(\y[0] ) );
    inv_1 \U1213/U907/U3  ( .x(\U1213/net4 ), .a(nbReset) );
    aoai211_1 \U1213/U1125/U28/U1/U1  ( .x(\U1213/U1125/U28/U1/clr ), .a(
        \U1213/nack[1] ), .b(\U1213/nack[0] ), .c(bsel), .d(nba) );
    nand3_1 \U1213/U1125/U28/U1/U2  ( .x(\U1213/U1125/U28/U1/set ), .a(bsel), 
        .b(\U1213/nack[1] ), .c(\U1213/nack[0] ) );
    nand2_2 \U1213/U1125/U28/U1/U3  ( .x(nba), .a(\U1213/U1125/U28/U1/clr ), 
        .b(\U1213/U1125/U28/U1/set ) );
    aoai211_1 \U1213/U1122/U28/U1/U1  ( .x(\U1213/U1122/U28/U1/clr ), .a(
        \U1213/nack[0] ), .b(\U1213/nack[1] ), .c(dsel), .d(nda) );
    nand3_1 \U1213/U1122/U28/U1/U2  ( .x(\U1213/U1122/U28/U1/set ), .a(dsel), 
        .b(\U1213/nack[0] ), .c(\U1213/nack[1] ) );
    nand2_2 \U1213/U1122/U28/U1/U3  ( .x(nda), .a(\U1213/U1122/U28/U1/clr ), 
        .b(\U1213/U1122/U28/U1/set ) );
    oa31_1 \U1213/U916_0_/U25/U1/Uclr  ( .x(\U1213/U916_0_/U25/U1/clr ), .a(
        nya), .b(\b[0] ), .c(\d[0] ), .d(\y[0] ) );
    oaoi211_1 \U1213/U916_0_/U25/U1/Uaoi  ( .x(\U1213/U916_0_/U25/U1/ob ), .a(
        \b[0] ), .b(\d[0] ), .c(nya), .d(\U1213/U916_0_/U25/U1/clr ) );
    inv_2 \U1213/U916_0_/U25/U1/Ui  ( .x(\y[0] ), .a(\U1213/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_1_/U25/U1/Uclr  ( .x(\U1213/U916_1_/U25/U1/clr ), .a(
        nya), .b(\b[1] ), .c(\d[1] ), .d(\y[1] ) );
    oaoi211_1 \U1213/U916_1_/U25/U1/Uaoi  ( .x(\U1213/U916_1_/U25/U1/ob ), .a(
        \b[1] ), .b(\d[1] ), .c(nya), .d(\U1213/U916_1_/U25/U1/clr ) );
    inv_2 \U1213/U916_1_/U25/U1/Ui  ( .x(\y[1] ), .a(\U1213/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_2_/U25/U1/Uclr  ( .x(\U1213/U916_2_/U25/U1/clr ), .a(
        nya), .b(\b[2] ), .c(\d[2] ), .d(\y[2] ) );
    oaoi211_1 \U1213/U916_2_/U25/U1/Uaoi  ( .x(\U1213/U916_2_/U25/U1/ob ), .a(
        \b[2] ), .b(\d[2] ), .c(nya), .d(\U1213/U916_2_/U25/U1/clr ) );
    inv_2 \U1213/U916_2_/U25/U1/Ui  ( .x(\y[2] ), .a(\U1213/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_3_/U25/U1/Uclr  ( .x(\U1213/U916_3_/U25/U1/clr ), .a(
        nya), .b(\b[3] ), .c(\d[3] ), .d(\y[3] ) );
    oaoi211_1 \U1213/U916_3_/U25/U1/Uaoi  ( .x(\U1213/U916_3_/U25/U1/ob ), .a(
        \b[3] ), .b(\d[3] ), .c(nya), .d(\U1213/U916_3_/U25/U1/clr ) );
    inv_2 \U1213/U916_3_/U25/U1/Ui  ( .x(\y[3] ), .a(\U1213/U916_3_/U25/U1/ob 
        ) );
    and3_2 \U1210/U1138/U9  ( .x(\d[3] ), .a(\cdh[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1137/U9  ( .x(\d[2] ), .a(\cdl[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1139/U9  ( .x(\d[1] ), .a(\cdh[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1210/U1136/U9  ( .x(\d[0] ), .a(\cdl[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1162/U1138/U9  ( .x(\a[3] ), .a(ih[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1137/U9  ( .x(\a[2] ), .a(il[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1139/U9  ( .x(\a[1] ), .a(ih[6]), .b(naa), .c(il[7]) );
    and3_2 \U1162/U1136/U9  ( .x(\a[0] ), .a(il[6]), .b(naa), .c(il[7]) );
    and3_2 \U1211/U1138/U9  ( .x(\b[3] ), .a(ih[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1137/U9  ( .x(\b[2] ), .a(il[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1139/U9  ( .x(\b[1] ), .a(ih[4]), .b(nba), .c(il[5]) );
    and3_2 \U1211/U1136/U9  ( .x(\b[0] ), .a(il[4]), .b(nba), .c(il[5]) );
    and3_2 \U1163/U1138/U9  ( .x(\c[3] ), .a(\cdh[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1137/U9  ( .x(\c[2] ), .a(\cdl[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1139/U9  ( .x(\c[1] ), .a(\cdh[2] ), .b(nca), .c(\cdl[3] )
         );
    and3_2 \U1163/U1136/U9  ( .x(\c[0] ), .a(\cdl[2] ), .b(nca), .c(\cdl[3] )
         );
    and2_1 \U1296/U1385/U8  ( .x(cg), .a(nbReset), .b(\U1296/ng ) );
    aoi222_1 \U1296/U1384/U30/U1  ( .x(\U1296/ng ), .a(nca), .b(net195), .c(
        nca), .d(\U1296/U1384/Z ), .e(net195), .f(\U1296/U1384/Z ) );
    inv_1 \U1296/U1384/U30/Uinv  ( .x(\U1296/U1384/Z ), .a(\U1296/ng ) );
    oa31_1 \U1296/U1386/U25/U1/Uclr  ( .x(\U1296/U1386/U25/U1/clr ), .a(
        \twobitack[2] ), .b(cg), .c(nca), .d(net195) );
    oaoi211_1 \U1296/U1386/U25/U1/Uaoi  ( .x(\U1296/U1386/U25/U1/ob ), .a(cg), 
        .b(nca), .c(\twobitack[2] ), .d(\U1296/U1386/U25/U1/clr ) );
    inv_2 \U1296/U1386/U25/U1/Ui  ( .x(net195), .a(\U1296/U1386/U25/U1/ob ) );
    and2_1 \U1298/U1385/U8  ( .x(dg), .a(nbReset), .b(\U1298/ng ) );
    aoi222_1 \U1298/U1384/U30/U1  ( .x(\U1298/ng ), .a(nda), .b(net193), .c(
        nda), .d(\U1298/U1384/Z ), .e(net193), .f(\U1298/U1384/Z ) );
    inv_1 \U1298/U1384/U30/Uinv  ( .x(\U1298/U1384/Z ), .a(\U1298/ng ) );
    oa31_1 \U1298/U1386/U25/U1/Uclr  ( .x(\U1298/U1386/U25/U1/clr ), .a(
        \twobitack[0] ), .b(dg), .c(nda), .d(net193) );
    oaoi211_1 \U1298/U1386/U25/U1/Uaoi  ( .x(\U1298/U1386/U25/U1/ob ), .a(dg), 
        .b(nda), .c(\twobitack[0] ), .d(\U1298/U1386/U25/U1/clr ) );
    inv_2 \U1298/U1386/U25/U1/Ui  ( .x(net193), .a(\U1298/U1386/U25/U1/ob ) );
    and2_1 \U1306/U1385/U8  ( .x(bg), .a(nbReset), .b(\U1306/ng ) );
    aoi222_1 \U1306/U1384/U30/U1  ( .x(\U1306/ng ), .a(nba), .b(\twobitack[1] 
        ), .c(nba), .d(\U1306/U1384/Z ), .e(\twobitack[1] ), .f(
        \U1306/U1384/Z ) );
    inv_1 \U1306/U1384/U30/Uinv  ( .x(\U1306/U1384/Z ), .a(\U1306/ng ) );
    oa31_1 \U1306/U1386/U25/U1/Uclr  ( .x(\U1306/U1386/U25/U1/clr ), .a(net199
        ), .b(bg), .c(nba), .d(\twobitack[1] ) );
    oaoi211_1 \U1306/U1386/U25/U1/Uaoi  ( .x(\U1306/U1386/U25/U1/ob ), .a(bg), 
        .b(nba), .c(net199), .d(\U1306/U1386/U25/U1/clr ) );
    inv_2 \U1306/U1386/U25/U1/Ui  ( .x(\twobitack[1] ), .a(
        \U1306/U1386/U25/U1/ob ) );
    and2_1 \U1295/U1385/U8  ( .x(ag), .a(nbReset), .b(\U1295/ng ) );
    aoi222_1 \U1295/U1384/U30/U1  ( .x(\U1295/ng ), .a(naa), .b(\twobitack[3] 
        ), .c(naa), .d(\U1295/U1384/Z ), .e(\twobitack[3] ), .f(
        \U1295/U1384/Z ) );
    inv_1 \U1295/U1384/U30/Uinv  ( .x(\U1295/U1384/Z ), .a(\U1295/ng ) );
    oa31_1 \U1295/U1386/U25/U1/Uclr  ( .x(\U1295/U1386/U25/U1/clr ), .a(net194
        ), .b(ag), .c(naa), .d(\twobitack[3] ) );
    oaoi211_1 \U1295/U1386/U25/U1/Uaoi  ( .x(\U1295/U1386/U25/U1/ob ), .a(ag), 
        .b(naa), .c(net194), .d(\U1295/U1386/U25/U1/clr ) );
    inv_2 \U1295/U1386/U25/U1/Ui  ( .x(\twobitack[3] ), .a(
        \U1295/U1386/U25/U1/ob ) );
    nand2_1 \U1297/U1131/U5  ( .x(\U1297/s ), .a(\U1297/r ), .b(\U1297/nback )
         );
    nand2_1 \U1297/U1103/U5  ( .x(\U1297/r ), .a(\U1297/naack ), .b(\U1297/s )
         );
    inv_1 \U1297/U1111/U3  ( .x(\U1297/reset ), .a(nbReset) );
    inv_1 \U1297/U1112/U3  ( .x(\U1297/naack ), .a(naa) );
    nor2_1 \U1297/U1130/U5  ( .x(\U1297/nback ), .a(nca), .b(\U1297/reset ) );
    aoai211_1 \U1297/U1128/U28/U1/U1  ( .x(\U1297/U1128/U28/U1/clr ), .a(
        \U1297/r ), .b(\U1297/naack ), .c(cg), .d(csel) );
    nand3_1 \U1297/U1128/U28/U1/U2  ( .x(\U1297/U1128/U28/U1/set ), .a(cg), 
        .b(\U1297/r ), .c(\U1297/naack ) );
    nand2_2 \U1297/U1128/U28/U1/U3  ( .x(csel), .a(\U1297/U1128/U28/U1/clr ), 
        .b(\U1297/U1128/U28/U1/set ) );
    aoai211_1 \U1297/U1127/U28/U1/U1  ( .x(\U1297/U1127/U28/U1/clr ), .a(
        \U1297/s ), .b(\U1297/nback ), .c(ag), .d(asel) );
    nand3_1 \U1297/U1127/U28/U1/U2  ( .x(\U1297/U1127/U28/U1/set ), .a(ag), 
        .b(\U1297/s ), .c(\U1297/nback ) );
    nand2_2 \U1297/U1127/U28/U1/U3  ( .x(asel), .a(\U1297/U1127/U28/U1/clr ), 
        .b(\U1297/U1127/U28/U1/set ) );
    nand2_1 \U1300/U1131/U5  ( .x(\U1300/s ), .a(\U1300/r ), .b(\U1300/nback )
         );
    nand2_1 \U1300/U1103/U5  ( .x(\U1300/r ), .a(\U1300/naack ), .b(\U1300/s )
         );
    inv_1 \U1300/U1111/U3  ( .x(\U1300/reset ), .a(nbReset) );
    inv_1 \U1300/U1112/U3  ( .x(\U1300/naack ), .a(nba) );
    nor2_1 \U1300/U1130/U5  ( .x(\U1300/nback ), .a(nda), .b(\U1300/reset ) );
    aoai211_1 \U1300/U1128/U28/U1/U1  ( .x(\U1300/U1128/U28/U1/clr ), .a(
        \U1300/r ), .b(\U1300/naack ), .c(dg), .d(dsel) );
    nand3_1 \U1300/U1128/U28/U1/U2  ( .x(\U1300/U1128/U28/U1/set ), .a(dg), 
        .b(\U1300/r ), .c(\U1300/naack ) );
    nand2_2 \U1300/U1128/U28/U1/U3  ( .x(dsel), .a(\U1300/U1128/U28/U1/clr ), 
        .b(\U1300/U1128/U28/U1/set ) );
    aoai211_1 \U1300/U1127/U28/U1/U1  ( .x(\U1300/U1127/U28/U1/clr ), .a(
        \U1300/s ), .b(\U1300/nback ), .c(bg), .d(bsel) );
    nand3_1 \U1300/U1127/U28/U1/U2  ( .x(\U1300/U1127/U28/U1/set ), .a(bg), 
        .b(\U1300/s ), .c(\U1300/nback ) );
    nand2_2 \U1300/U1127/U28/U1/U3  ( .x(bsel), .a(\U1300/U1127/U28/U1/clr ), 
        .b(\U1300/U1127/U28/U1/set ) );
    aoai211_1 \U1289/U1150/U28/U1/U1  ( .x(\U1289/U1150/U28/U1/clr ), .a(il[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[2] ) );
    nand3_1 \U1289/U1150/U28/U1/U2  ( .x(\U1289/U1150/U28/U1/set ), .a(net195), 
        .b(il[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1150/U28/U1/U3  ( .x(\cdl[2] ), .a(
        \U1289/U1150/U28/U1/clr ), .b(\U1289/U1150/U28/U1/set ) );
    aoai211_1 \U1289/U1152/U28/U1/U1  ( .x(\U1289/U1152/U28/U1/clr ), .a(il[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[3] ) );
    nand3_1 \U1289/U1152/U28/U1/U2  ( .x(\U1289/U1152/U28/U1/set ), .a(net195), 
        .b(il[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1152/U28/U1/U3  ( .x(\cdl[3] ), .a(
        \U1289/U1152/U28/U1/clr ), .b(\U1289/U1152/U28/U1/set ) );
    aoai211_1 \U1289/U1149/U28/U1/U1  ( .x(\U1289/U1149/U28/U1/clr ), .a(ih[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[2] ) );
    nand3_1 \U1289/U1149/U28/U1/U2  ( .x(\U1289/U1149/U28/U1/set ), .a(net195), 
        .b(ih[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1149/U28/U1/U3  ( .x(\cdh[2] ), .a(
        \U1289/U1149/U28/U1/clr ), .b(\U1289/U1149/U28/U1/set ) );
    aoai211_1 \U1289/U1151/U28/U1/U1  ( .x(\U1289/U1151/U28/U1/clr ), .a(ih[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[3] ) );
    nand3_1 \U1289/U1151/U28/U1/U2  ( .x(\U1289/U1151/U28/U1/set ), .a(net195), 
        .b(ih[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1151/U28/U1/U3  ( .x(\cdh[3] ), .a(
        \U1289/U1151/U28/U1/clr ), .b(\U1289/U1151/U28/U1/set ) );
    inv_1 \U1289/U1148/U1147/U3  ( .x(\U1289/U1148/net189 ), .a(
        \U1289/bnreset ) );
    nor2_1 \U1289/U1148/U582/U5  ( .x(\U1289/U1148/net192 ), .a(\cdl[3] ), .b(
        \cdh[3] ) );
    nor2_1 \U1289/U1148/U580/U5  ( .x(\U1289/U1148/net191 ), .a(\cdl[2] ), .b(
        \cdh[2] ) );
    nor2_2 \U1289/U1148/U1146/U6  ( .x(\twobitack[2] ), .a(
        \U1289/U1148/net190 ), .b(\U1289/U1148/net189 ) );
    aoi222_1 \U1289/U1148/U1141/U30/U1  ( .x(\U1289/U1148/net190 ), .a(
        \U1289/U1148/net191 ), .b(\U1289/U1148/net192 ), .c(
        \U1289/U1148/net191 ), .d(\U1289/U1148/U1141/Z ), .e(
        \U1289/U1148/net192 ), .f(\U1289/U1148/U1141/Z ) );
    inv_1 \U1289/U1148/U1141/U30/Uinv  ( .x(\U1289/U1148/U1141/Z ), .a(
        \U1289/U1148/net190 ) );
    aoai211_1 \U1271/U1150/U28/U1/U1  ( .x(\U1271/U1150/U28/U1/clr ), .a(il[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[0] ) );
    nand3_1 \U1271/U1150/U28/U1/U2  ( .x(\U1271/U1150/U28/U1/set ), .a(net193), 
        .b(il[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1150/U28/U1/U3  ( .x(\cdl[0] ), .a(
        \U1271/U1150/U28/U1/clr ), .b(\U1271/U1150/U28/U1/set ) );
    aoai211_1 \U1271/U1152/U28/U1/U1  ( .x(\U1271/U1152/U28/U1/clr ), .a(il[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[1] ) );
    nand3_1 \U1271/U1152/U28/U1/U2  ( .x(\U1271/U1152/U28/U1/set ), .a(net193), 
        .b(il[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1152/U28/U1/U3  ( .x(\cdl[1] ), .a(
        \U1271/U1152/U28/U1/clr ), .b(\U1271/U1152/U28/U1/set ) );
    aoai211_1 \U1271/U1149/U28/U1/U1  ( .x(\U1271/U1149/U28/U1/clr ), .a(ih[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[0] ) );
    nand3_1 \U1271/U1149/U28/U1/U2  ( .x(\U1271/U1149/U28/U1/set ), .a(net193), 
        .b(ih[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1149/U28/U1/U3  ( .x(\cdh[0] ), .a(
        \U1271/U1149/U28/U1/clr ), .b(\U1271/U1149/U28/U1/set ) );
    aoai211_1 \U1271/U1151/U28/U1/U1  ( .x(\U1271/U1151/U28/U1/clr ), .a(ih[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[1] ) );
    nand3_1 \U1271/U1151/U28/U1/U2  ( .x(\U1271/U1151/U28/U1/set ), .a(net193), 
        .b(ih[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1151/U28/U1/U3  ( .x(\cdh[1] ), .a(
        \U1271/U1151/U28/U1/clr ), .b(\U1271/U1151/U28/U1/set ) );
    inv_1 \U1271/U1148/U1147/U3  ( .x(\U1271/U1148/net189 ), .a(
        \U1271/bnreset ) );
    nor2_1 \U1271/U1148/U582/U5  ( .x(\U1271/U1148/net192 ), .a(\cdl[1] ), .b(
        \cdh[1] ) );
    nor2_1 \U1271/U1148/U580/U5  ( .x(\U1271/U1148/net191 ), .a(\cdl[0] ), .b(
        \cdh[0] ) );
    nor2_2 \U1271/U1148/U1146/U6  ( .x(\twobitack[0] ), .a(
        \U1271/U1148/net190 ), .b(\U1271/U1148/net189 ) );
    aoi222_1 \U1271/U1148/U1141/U30/U1  ( .x(\U1271/U1148/net190 ), .a(
        \U1271/U1148/net191 ), .b(\U1271/U1148/net192 ), .c(
        \U1271/U1148/net191 ), .d(\U1271/U1148/U1141/Z ), .e(
        \U1271/U1148/net192 ), .f(\U1271/U1148/U1141/Z ) );
    inv_1 \U1271/U1148/U1141/U30/Uinv  ( .x(\U1271/U1148/U1141/Z ), .a(
        \U1271/U1148/net190 ) );
    nand2_1 \U1225/U1128/U5  ( .x(\U1225/s ), .a(\U1225/r ), .b(\U1225/nback )
         );
    nand2_1 \U1225/U1103/U5  ( .x(\U1225/r ), .a(\U1225/naack ), .b(\U1225/s )
         );
    inv_1 \U1225/U1111/U3  ( .x(\U1225/reset ), .a(nbReset) );
    inv_1 \U1225/U1112/U3  ( .x(\U1225/naack ), .a(nxa) );
    nor2_1 \U1225/U1127/U5  ( .x(\U1225/nback ), .a(nyla), .b(\U1225/reset )
         );
    and2_2 \U1225/U1129/U8  ( .x(xsel), .a(\U1225/nback ), .b(\U1225/s ) );
    and2_2 \U1225/U1124/U8  ( .x(ysel), .a(\U1225/r ), .b(\U1225/naack ) );
    and3_4 \U1308/U20/U9  ( .x(nya), .a(\U1308/nack[1] ), .b(\U1308/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U1308/U18/U5  ( .x(\U1308/nack[0] ), .a(\yl[3] ), .b(\yl[0] ) );
    nor2_1 \U1308/U19/U5  ( .x(\U1308/nack[1] ), .a(\yl[1] ), .b(\yl[2] ) );
    ao222_2 \U1308/U15_0_/U19/U1/U1  ( .x(\yl[0] ), .a(\y[0] ), .b(nyla), .c(
        \y[0] ), .d(\yl[0] ), .e(nyla), .f(\yl[0] ) );
    ao222_2 \U1308/U15_1_/U19/U1/U1  ( .x(\yl[1] ), .a(\y[1] ), .b(nyla), .c(
        \y[1] ), .d(\yl[1] ), .e(nyla), .f(\yl[1] ) );
    ao222_2 \U1308/U15_2_/U19/U1/U1  ( .x(\yl[2] ), .a(\y[2] ), .b(nyla), .c(
        \y[2] ), .d(\yl[2] ), .e(nyla), .f(\yl[2] ) );
    ao222_2 \U1308/U15_3_/U19/U1/U1  ( .x(\yl[3] ), .a(\y[3] ), .b(nyla), .c(
        \y[3] ), .d(\yl[3] ), .e(nyla), .f(\yl[3] ) );
    buf_3 U1 ( .x(\U1271/bnreset ), .a(nbReset) );
    buf_3 U2 ( .x(\U1289/bnreset ), .a(nbReset) );
endmodule


module chain_dr8bit_completion_44 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_45 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_46 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_47 ( o, i );
input  [15:0] i;
output o;
    wire y, \ny[3] , \ny[2] , \ny[1] , \ny[0] , x, \nx[3] , \nx[2] , \nx[1] , 
        \nx[0] , \U6/Z , \U3/net2 , \U3/net3 , \U3/U20/Z , \U3/U21/Z , 
        \U3/U19/Z , \U5/net2 , \U5/net3 , \U5/U20/Z , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr32bit_completion_10 ( o, i );
input  [63:0] i;
output o;
    wire nx, \cd[3] , \cd[2] , ny, \cd[0] , \cd[1] , \U16/Z , \U6/Z , \U15/Z ;
    chain_dr8bit_completion_44 U11 ( .o(\cd[3] ), .i({i[63], i[62], i[61], 
        i[60], i[59], i[58], i[57], i[56], i[31], i[30], i[29], i[28], i[27], 
        i[26], i[25], i[24]}) );
    chain_dr8bit_completion_47 U14 ( .o(\cd[2] ), .i({i[55], i[54], i[53], 
        i[52], i[51], i[50], i[49], i[48], i[23], i[22], i[21], i[20], i[19], 
        i[18], i[17], i[16]}) );
    chain_dr8bit_completion_46 U13 ( .o(\cd[1] ), .i({i[47], i[46], i[45], 
        i[44], i[43], i[42], i[41], i[40], i[15], i[14], i[13], i[12], i[11], 
        i[10], i[9], i[8]}) );
    chain_dr8bit_completion_45 U12 ( .o(\cd[0] ), .i({i[39], i[38], i[37], 
        i[36], i[35], i[34], i[33], i[32], i[7], i[6], i[5], i[4], i[3], i[2], 
        i[1], i[0]}) );
    aoi222_1 \U16/U30/U1  ( .x(ny), .a(\cd[0] ), .b(\cd[1] ), .c(\cd[0] ), .d(
        \U16/Z ), .e(\cd[1] ), .f(\U16/Z ) );
    inv_1 \U16/U30/Uinv  ( .x(\U16/Z ), .a(ny) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(ny), .b(nx), .c(ny), .d(\U6/Z ), .e(nx), 
        .f(\U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U15/U30/U1  ( .x(nx), .a(\cd[3] ), .b(\cd[2] ), .c(\cd[3] ), .d(
        \U15/Z ), .e(\cd[2] ), .f(\U15/Z ) );
    inv_1 \U15/U30/Uinv  ( .x(\U15/Z ), .a(nx) );
endmodule


module chain_selement_ga_72 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_73 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_t_ctrl_2 ( cack, fcdefer, fcslowack, screq, ack, defer, fcack, 
    nReset, scack, slowack );
input  ack, defer, fcack, nReset, scack, slowack;
output cack, fcdefer, fcslowack, screq;
    wire net269, net280, net275, net270, net265, net278, net276, net277, 
        net263, net271, net266, net279, net272, net264, net267, net273, net268, 
        net274, \U49/U28/U1/clr , \U49/U28/U1/set , \U50/U28/U1/clr , 
        \U50/U28/U1/set , \U51/U28/U1/clr , \U51/U28/U1/set , \U57/acb , 
        \U57/U1/Z ;
    chain_selement_ga_73 U55 ( .Aa(net269), .Br(fcdefer), .Ar(net280), .Ba(
        fcack) );
    chain_selement_ga_72 U54 ( .Aa(net275), .Br(fcslowack), .Ar(net270), .Ba(
        fcack) );
    or2_4 \U12/U12  ( .x(net268), .a(net266), .b(net270) );
    or2_4 \U56/U12  ( .x(net274), .a(net275), .b(net269) );
    or2_4 \U14/U12  ( .x(net273), .a(net274), .b(net266) );
    or3_1 \U36/U12  ( .x(cack), .a(net267), .b(net264), .c(net272) );
    nor3_1 \U21/U7  ( .x(net271), .a(net270), .b(net266), .c(net280) );
    and2_1 \U53/U8  ( .x(net263), .a(net271), .b(nReset) );
    and2_1 \U43/U8  ( .x(net277), .a(net265), .b(nReset) );
    nor2_1 \U22/U5  ( .x(net265), .a(net278), .b(net276) );
    ao222_2 \U44/U19/U1/U1  ( .x(net276), .a(net280), .b(net273), .c(net280), 
        .d(net276), .e(net273), .f(net276) );
    ao222_2 \U40/U19/U1/U1  ( .x(net280), .a(net272), .b(net277), .c(net272), 
        .d(net280), .e(net277), .f(net280) );
    ao222_2 \U45/U19/U1/U1  ( .x(net279), .a(net273), .b(net268), .c(net273), 
        .d(net279), .e(net268), .f(net279) );
    ao222_2 \U42/U19/U1/U1  ( .x(net266), .a(net277), .b(net267), .c(net277), 
        .d(net266), .e(net267), .f(net266) );
    ao222_2 \U39/U19/U1/U1  ( .x(net270), .a(net277), .b(net264), .c(net277), 
        .d(net270), .e(net264), .f(net270) );
    aoai211_1 \U49/U28/U1/U1  ( .x(\U49/U28/U1/clr ), .a(ack), .b(nReset), .c(
        net263), .d(net267) );
    nand3_1 \U49/U28/U1/U2  ( .x(\U49/U28/U1/set ), .a(net263), .b(ack), .c(
        nReset) );
    nand2_2 \U49/U28/U1/U3  ( .x(net267), .a(\U49/U28/U1/clr ), .b(
        \U49/U28/U1/set ) );
    aoai211_1 \U50/U28/U1/U1  ( .x(\U50/U28/U1/clr ), .a(slowack), .b(nReset), 
        .c(net263), .d(net264) );
    nand3_1 \U50/U28/U1/U2  ( .x(\U50/U28/U1/set ), .a(net263), .b(slowack), 
        .c(nReset) );
    nand2_2 \U50/U28/U1/U3  ( .x(net264), .a(\U50/U28/U1/clr ), .b(
        \U50/U28/U1/set ) );
    aoai211_1 \U51/U28/U1/U1  ( .x(\U51/U28/U1/clr ), .a(defer), .b(nReset), 
        .c(net263), .d(net272) );
    nand2_2 \U51/U28/U1/U3  ( .x(net272), .a(\U51/U28/U1/clr ), .b(
        \U51/U28/U1/set ) );
    and2_1 \U57/U2/U8  ( .x(screq), .a(net279), .b(\U57/acb ) );
    nor2_1 \U57/U3/U5  ( .x(net278), .a(\U57/acb ), .b(scack) );
    oai21_1 \U57/U1/U30/U1/U1  ( .x(\U57/acb ), .a(\U57/U1/Z ), .b(scack), .c(
        net279) );
    inv_1 \U57/U1/U30/U1/U2  ( .x(\U57/U1/Z ), .a(\U57/acb ) );
    nand3_0 U1 ( .x(\U51/U28/U1/set ), .a(net263), .b(defer), .c(nReset) );
endmodule


module chain_mergepackets_5 ( naa, nba, o, a, b, nReset, noa );
output [4:0] o;
input  [4:0] a;
input  [4:0] b;
input  nReset, noa;
output naa, nba;
    wire \noack[1] , \noack[0] , reset, bsel, as, setb, asel, seta, 
        \U916_0_/U25/U1/clr , \U916_0_/U25/U1/ob , \U916_1_/U25/U1/clr , 
        \U916_1_/U25/U1/ob , \U916_2_/U25/U1/clr , \U916_2_/U25/U1/ob , 
        \U916_3_/U25/U1/clr , \U916_3_/U25/U1/ob ;
    and2_1 \U1155/U8  ( .x(as), .a(seta), .b(asel) );
    nand2_1 \U1145/U5  ( .x(asel), .a(bsel), .b(seta) );
    nand2_1 \U1103/U5  ( .x(bsel), .a(setb), .b(asel) );
    inv_1 \U1135/U3  ( .x(reset), .a(nReset) );
    inv_1 \U1134/U3  ( .x(setb), .a(a[4]) );
    and3_2 \U1154/U9  ( .x(naa), .a(\noack[1] ), .b(\noack[0] ), .c(as) );
    nor3_1 \U1127/U7  ( .x(\noack[0] ), .a(o[1]), .b(reset), .c(o[0]) );
    nor2_1 \U1132/U5  ( .x(\noack[1] ), .a(o[3]), .b(o[2]) );
    oa31_1 \U916_0_/U25/U1/Uclr  ( .x(\U916_0_/U25/U1/clr ), .a(noa), .b(a[0]), 
        .c(b[0]), .d(o[0]) );
    oaoi211_1 \U916_0_/U25/U1/Uaoi  ( .x(\U916_0_/U25/U1/ob ), .a(a[0]), .b(b
        [0]), .c(noa), .d(\U916_0_/U25/U1/clr ) );
    inv_2 \U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U916_0_/U25/U1/ob ) );
    oa31_1 \U916_1_/U25/U1/Uclr  ( .x(\U916_1_/U25/U1/clr ), .a(noa), .b(a[1]), 
        .c(b[1]), .d(o[1]) );
    oaoi211_1 \U916_1_/U25/U1/Uaoi  ( .x(\U916_1_/U25/U1/ob ), .a(a[1]), .b(b
        [1]), .c(noa), .d(\U916_1_/U25/U1/clr ) );
    inv_2 \U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U916_1_/U25/U1/ob ) );
    oa31_1 \U916_2_/U25/U1/Uclr  ( .x(\U916_2_/U25/U1/clr ), .a(noa), .b(a[2]), 
        .c(b[2]), .d(o[2]) );
    oaoi211_1 \U916_2_/U25/U1/Uaoi  ( .x(\U916_2_/U25/U1/ob ), .a(a[2]), .b(b
        [2]), .c(noa), .d(\U916_2_/U25/U1/clr ) );
    inv_2 \U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U916_2_/U25/U1/ob ) );
    oa31_1 \U916_3_/U25/U1/Uclr  ( .x(\U916_3_/U25/U1/clr ), .a(noa), .b(a[3]), 
        .c(b[3]), .d(o[3]) );
    oaoi211_1 \U916_3_/U25/U1/Uaoi  ( .x(\U916_3_/U25/U1/ob ), .a(a[3]), .b(b
        [3]), .c(noa), .d(\U916_3_/U25/U1/clr ) );
    inv_2 \U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U916_3_/U25/U1/ob ) );
    ao222_2 \U1148/U19/U1/U1  ( .x(o[4]), .a(noa), .b(b[4]), .c(noa), .d(o[4]), 
        .e(b[4]), .f(o[4]) );
    aoi21_1 \U1153/U11  ( .x(seta), .a(o[4]), .b(setb), .c(reset) );
    and3_3 U1 ( .x(nba), .a(bsel), .b(\noack[0] ), .c(\noack[1] ) );
endmodule


module target_dmem ( addr, ccol, chainresponse, crnw, csize, ctag, lock, 
    nchaincommandack, nrouteack, pred, rack, routetxreq, seq, tag_h, tag_l, wd, 
    cack, cdefer, chaincommand, cndefer, cok, err, nReset, nchainresponseack, 
    rd, route, routetxack );
output [63:0] addr;
output [5:0] ccol;
output [4:0] chainresponse;
output [1:0] crnw;
output [3:0] csize;
output [9:0] ctag;
output [1:0] lock;
output [1:0] pred;
output [1:0] seq;
output [4:0] tag_h;
output [4:0] tag_l;
output [63:0] wd;
input  [4:0] chaincommand;
input  [1:0] err;
input  [63:0] rd;
input  [4:0] route;
input  cack, cdefer, cndefer, cok, nReset, nchainresponseack, routetxack;
output nchaincommandack, nrouteack, rack, routetxreq;
    wire n10, n11, n12, n13, n14, \net242[0] , \net242[1] , \net242[2] , 
        \net242[3] , \net242[4] , \net242[5] , \net242[6] , \net242[7] , 
        \net242[8] , \net242[9] , \net242[10] , \net243[0] , \net243[1] , 
        \net243[2] , \net243[3] , \net243[4] , \net243[5] , \net243[6] , 
        \net243[7] , \net243[8] , \net243[9] , \net243[10] , \net244[0] , 
        \net244[1] , \net244[2] , \net244[3] , \net244[4] , \net244[5] , 
        \net244[6] , \net244[7] , \net244[8] , \net244[9] , \net244[10] , 
        \chainff_l[7] , \chainff_l[6] , \chainff_l[5] , \chainff_l[4] , 
        \chainff_l[3] , \chainff_l[2] , \chainff_l[1] , \chainff_l[0] , 
        \chdrack[0] , \chdrack[1] , \obl[7] , \obl[6] , \obl[5] , \obl[4] , 
        \obl[3] , \obl[2] , \obl[1] , \obl[0] , \tcbh[7] , \tcbh[6] , 
        \tcbh[5] , \tcbh[4] , \tcbh[3] , \tcbh[2] , \tcbh[1] , \tcbh[0] , 
        \tcbl[7] , \tcbl[6] , \tcbl[5] , \tcbl[4] , \tcbl[3] , \tcbl[2] , 
        \tcbl[1] , \tcbl[0] , \tresponse[4] , \tresponse[3] , \tresponse[2] , 
        \tresponse[1] , \tresponse[0] , \nchdr_ack[10] , \nchdr_ack[9] , 
        \nchdr_ack[8] , \nchdr_ack[7] , \nchdr_ack[6] , \nchdr_ack[5] , 
        \nchdr_ack[4] , \nchdr_ack[3] , \nchdr_ack[2] , \nchdr_ack[1] , 
        \nchdr_ack[0] , \chainff_h[7] , \chainff_h[6] , \chainff_h[5] , 
        \chainff_h[4] , \chainff_h[3] , \chainff_h[2] , \chainff_h[1] , 
        \chainff_h[0] , \rhdr_l[15] , \rhdr_l[14] , \rhdr_l[13] , \rhdr_l[7] , 
        \rhdr_l[6] , \rhdr_l[5] , \obh[7] , \obh[6] , \obh[5] , \obh[4] , 
        \obh[3] , \obh[2] , \obh[1] , \obh[0] , \rhdr_h[15] , \rhdr_h[14] , 
        \rhdr_h[13] , \rhdr_h[7] , \rhdr_h[6] , \rhdr_h[5] , net265, nbreset, 
        net248, rhdrack, read_ctrlack, chainff_ack, read_req, read_cd, teop, 
        fcack, tcba, net145, screq, fcslowack, fcdefer, read_ack, 
        ntresponseack, net200, noba, pullcd, net168, net188, net201, net194, 
        net178, net189, net191, net284, hdrcd, chdrctrlack, \U1770/U21/nr , 
        \U1770/U21/nd , \U1770/U21/n2 , \U1761/U28/Z , \U1761/U32/Z , 
        \U1761/U29/Z , \U1761/U33/Z , \U1761/U30/Z , \U1761/U31/Z , \U1632/Z , 
        \U1676/Z , \U1761/y[0] , \U1761/y[1] , \U1761/x[1] , \U1761/x[3] , 
        \U1761/x[2] , \U1761/x[0] , \U1574_0_/net231 , \U1574_1_/net231 , 
        \U1574_2_/net231 , \U1574_3_/net231 , \U1574_4_/net231 , 
        \U1574_5_/net231 , \U1574_6_/net231 , \U1574_7_/net231 , 
        \U1574_8_/net231 , \U1574_9_/net231 , \U1574_10_/net231 , n6, n7, n8, 
        n9;
    chain_sendword_2 U1765 ( .ctrlack(read_ctrlack), .oh({\chainff_h[7] , 
        \chainff_h[6] , \chainff_h[5] , \chainff_h[4] , \chainff_h[3] , 
        \chainff_h[2] , \chainff_h[1] , \chainff_h[0] }), .ol({\chainff_l[7] , 
        \chainff_l[6] , \chainff_l[5] , \chainff_l[4] , \chainff_l[3] , 
        \chainff_l[2] , \chainff_l[1] , \chainff_l[0] }), .chainackff(
        chainff_ack), .ctrlreq(read_req), .ih(rd[63:32]), .il(rd[31:0]) );
    chain_dr32bit_completion_10 rd_cd ( .o(read_cd), .i(rd) );
    chain_trhdr_2 xmitHdr ( .chainff_ack(chainff_ack), .chainh({\tcbh[7] , 
        \tcbh[6] , \tcbh[5] , \tcbh[4] , \tcbh[3] , \tcbh[2] , \tcbh[1] , 
        \tcbh[0] }), .chainl({\tcbl[7] , \tcbl[6] , \tcbl[5] , \tcbl[4] , 
        \tcbl[3] , \tcbl[2] , \tcbl[1] , \tcbl[0] }), .eop(teop), .hdrack(
        rhdrack), .normal_ack(rack), .notify_ack(fcack), .read_req(read_req), 
        .routereq(routetxreq), .chain_ff_h({\chainff_h[7] , \chainff_h[6] , 
        \chainff_h[5] , \chainff_h[4] , \chainff_h[3] , \chainff_h[2] , 
        \chainff_h[1] , \chainff_h[0] }), .chainack(tcba), .chainff_l({
        \chainff_l[7] , \chainff_l[6] , \chainff_l[5] , \chainff_l[4] , 
        \chainff_l[3] , \chainff_l[2] , \chainff_l[1] , \chainff_l[0] }), 
        .eopack(net145), .err(err), .nReset(n6), .normal_response(screq), 
        .notify_accept(fcslowack), .notify_defer(fcdefer), .rcol_h({
        \rhdr_h[15] , \rhdr_h[14] , \rhdr_h[13] }), .rcol_l({\rhdr_l[15] , 
        \rhdr_l[14] , \rhdr_l[13] }), .read_ack(read_ack), .rnw_h(\rhdr_h[7] ), 
        .rnw_l(\rhdr_l[7] ), .routeack(routetxack), .rsize_h({\rhdr_h[6] , 
        \rhdr_h[5] }), .rsize_l({\rhdr_l[6] , \rhdr_l[5] }), .rtag_h(tag_h), 
        .rtag_l(tag_l) );
    chain_dr2fr_byte_5 dr2fr ( .eop_ack(net145), .ia(tcba), .o({\tresponse[4] , 
        \tresponse[3] , \tresponse[2] , \tresponse[1] , \tresponse[0] }), 
        .eop(teop), .ih({\tcbh[7] , \tcbh[6] , \tcbh[5] , \tcbh[4] , \tcbh[3] , 
        \tcbh[2] , \tcbh[1] , \tcbh[0] }), .il({\tcbl[7] , \tcbl[6] , 
        \tcbl[5] , \tcbl[4] , \tcbl[3] , \tcbl[2] , \tcbl[1] , \tcbl[0] }), 
        .nReset(nbreset), .noa(ntresponseack) );
    chain_mergepackets_5 merger ( .naa(nrouteack), .nba(ntresponseack), .o(
        chainresponse), .a(route), .b({\tresponse[4] , \tresponse[3] , 
        \tresponse[2] , \tresponse[1] , \tresponse[0] }), .nReset(nbreset), 
        .noa(nchainresponseack) );
    chain_tchdr_2 header ( .addr_req(net200), .col_h(ccol[5:3]), .col_l(ccol
        [2:0]), .itag_h(ctag[9:5]), .itag_l(ctag[4:0]), .lock(lock), .ncback(
        noba), .pred(pred), .pullcd(pullcd), .reset(net168), .rnw_h(n10), 
        .rnw_l(n11), .seq(seq), .size_h({n12, csize[2]}), .size_l({n13, n14}), 
        .write_req(net188), .chwh({\obh[7] , \obh[6] , \obh[5] , \obh[4] , 
        \obh[3] , \obh[2] , \obh[1] , \obh[0] }), .chwl({\obl[7] , \obl[6] , 
        \obl[5] , \obl[4] , \obl[3] , \obl[2] , \obl[1] , \obl[0] }), 
        .addr_ack(net201), .addr_pull(net194), .nReset(n6), .nack(net178), 
        .write_ack(net189), .write_pull(net191) );
    chain_irdemux_32new_5 wd_hld ( .ctrlack(net189), .oh(wd[63:32]), .ol(wd
        [31:0]), .pullreq(net191), .pull_h({\obh[7] , \obh[6] , \obh[5] , 
        \obh[4] , \obh[3] , \obh[2] , \obh[1] , \obh[0] }), .pull_l({\obl[7] , 
        \obl[6] , \obl[5] , \obl[4] , \obl[3] , \obl[2] , \obl[1] , \obl[0] }), 
        .pullcd(pullcd), .reset(net168), .ctrlreq(net188) );
    chain_irdemux_32new_4 adr_hld ( .ctrlack(net201), .oh(addr[63:32]), .ol(
        addr[31:0]), .pullreq(net194), .pull_h({\obh[7] , \obh[6] , \obh[5] , 
        \obh[4] , \obh[3] , \obh[2] , \obh[1] , \obh[0] }), .pull_l({\obl[7] , 
        \obl[6] , \obl[5] , \obl[4] , \obl[3] , \obl[2] , \obl[1] , \obl[0] }), 
        .pullcd(pullcd), .reset(net168), .ctrlreq(net200) );
    chain_fr2dr_byte_2 chain_decoder ( .nia(nchaincommandack), .oh({\obh[7] , 
        \obh[6] , \obh[5] , \obh[4] , \obh[3] , \obh[2] , \obh[1] , \obh[0] }), 
        .ol({\obl[7] , \obl[6] , \obl[5] , \obl[4] , \obl[3] , \obl[2] , 
        \obl[1] , \obl[0] }), .i(chaincommand), .nReset(nbreset), .noa(noba)
         );
    chain_t_ctrl_2 cmd_ctrl ( .cack(net284), .fcdefer(fcdefer), .fcslowack(
        fcslowack), .screq(screq), .ack(cok), .defer(cdefer), .fcack(fcack), 
        .nReset(n6), .scack(rack), .slowack(cndefer) );
    inv_1 \I4/U3  ( .x(net265), .a(nbreset) );
    ao222_1 \U1761/U37/U18/U1/U1  ( .x(\chdrack[0] ), .a(\U1761/y[0] ), .b(
        \U1761/y[1] ), .c(\U1761/y[0] ), .d(\chdrack[0] ), .e(\U1761/y[1] ), 
        .f(\chdrack[0] ) );
    ao222_1 \U1762/U18/U1/U1  ( .x(chdrctrlack), .a(hdrcd), .b(net284), .c(
        hdrcd), .d(chdrctrlack), .e(net284), .f(chdrctrlack) );
    ao222_1 \U1769/U18/U1/U1  ( .x(read_ack), .a(read_ctrlack), .b(read_cd), 
        .c(read_ctrlack), .d(read_ack), .e(read_cd), .f(read_ack) );
    aoi222_1 \U1761/U28/U30/U1  ( .x(\U1761/x[3] ), .a(\nchdr_ack[7] ), .b(
        \nchdr_ack[6] ), .c(\nchdr_ack[7] ), .d(\U1761/U28/Z ), .e(
        \nchdr_ack[6] ), .f(\U1761/U28/Z ) );
    inv_1 \U1761/U28/U30/Uinv  ( .x(\U1761/U28/Z ), .a(\U1761/x[3] ) );
    aoi222_1 \U1761/U32/U30/U1  ( .x(\U1761/x[0] ), .a(\nchdr_ack[1] ), .b(
        \nchdr_ack[0] ), .c(\nchdr_ack[1] ), .d(\U1761/U32/Z ), .e(
        \nchdr_ack[0] ), .f(\U1761/U32/Z ) );
    inv_1 \U1761/U32/U30/Uinv  ( .x(\U1761/U32/Z ), .a(\U1761/x[0] ) );
    aoi222_1 \U1761/U29/U30/U1  ( .x(\U1761/x[2] ), .a(\nchdr_ack[5] ), .b(
        \nchdr_ack[4] ), .c(\nchdr_ack[5] ), .d(\U1761/U29/Z ), .e(
        \nchdr_ack[4] ), .f(\U1761/U29/Z ) );
    inv_1 \U1761/U29/U30/Uinv  ( .x(\U1761/U29/Z ), .a(\U1761/x[2] ) );
    aoi222_1 \U1761/U33/U30/U1  ( .x(\U1761/y[0] ), .a(\U1761/x[1] ), .b(
        \U1761/x[0] ), .c(\U1761/x[1] ), .d(\U1761/U33/Z ), .e(\U1761/x[0] ), 
        .f(\U1761/U33/Z ) );
    inv_1 \U1761/U33/U30/Uinv  ( .x(\U1761/U33/Z ), .a(\U1761/y[0] ) );
    aoi222_1 \U1761/U30/U30/U1  ( .x(\U1761/y[1] ), .a(\U1761/x[3] ), .b(
        \U1761/x[2] ), .c(\U1761/x[3] ), .d(\U1761/U30/Z ), .e(\U1761/x[2] ), 
        .f(\U1761/U30/Z ) );
    inv_1 \U1761/U30/U30/Uinv  ( .x(\U1761/U30/Z ), .a(\U1761/y[1] ) );
    aoi222_1 \U1761/U31/U30/U1  ( .x(\U1761/x[1] ), .a(\nchdr_ack[3] ), .b(
        \nchdr_ack[2] ), .c(\nchdr_ack[3] ), .d(\U1761/U31/Z ), .e(
        \nchdr_ack[2] ), .f(\U1761/U31/Z ) );
    inv_1 \U1761/U31/U30/Uinv  ( .x(\U1761/U31/Z ), .a(\U1761/x[1] ) );
    aoi222_1 \U1632/U30/U1  ( .x(net178), .a(cack), .b(chdrctrlack), .c(cack), 
        .d(\U1632/Z ), .e(chdrctrlack), .f(\U1632/Z ) );
    inv_1 \U1632/U30/Uinv  ( .x(\U1632/Z ), .a(net178) );
    aoi222_1 \U1676/U30/U1  ( .x(hdrcd), .a(\chdrack[0] ), .b(\chdrack[1] ), 
        .c(\chdrack[0] ), .d(\U1676/Z ), .e(\chdrack[1] ), .f(\U1676/Z ) );
    inv_1 \U1676/U30/Uinv  ( .x(\U1676/Z ), .a(hdrcd) );
    nor3_1 \U1770/U21/Unr  ( .x(\U1770/U21/nr ), .a(\nchdr_ack[10] ), .b(
        \nchdr_ack[9] ), .c(\nchdr_ack[8] ) );
    nand3_1 \U1770/U21/Und  ( .x(\U1770/U21/nd ), .a(\nchdr_ack[10] ), .b(
        \nchdr_ack[9] ), .c(\nchdr_ack[8] ) );
    oa21_1 \U1770/U21/U1  ( .x(\U1770/U21/n2 ), .a(\U1770/U21/n2 ), .b(
        \U1770/U21/nr ), .c(\U1770/U21/nd ) );
    inv_1 \U1770/U21/U3  ( .x(\chdrack[1] ), .a(\U1770/U21/n2 ) );
    nor2_1 \U1652_0_/U2/U5  ( .x(\nchdr_ack[0] ), .a(\net242[10] ), .b(
        \net244[10] ) );
    ao222_2 \U1652_0_/U12/U19/U1/U1  ( .x(\net244[10] ), .a(\net243[10] ), .b(
        csize[0]), .c(\net243[10] ), .d(\net244[10] ), .e(csize[0]), .f(
        \net244[10] ) );
    ao222_2 \U1652_0_/U11/U19/U1/U1  ( .x(\net242[10] ), .a(csize[2]), .b(
        \net243[10] ), .c(csize[2]), .d(\net242[10] ), .e(\net243[10] ), .f(
        \net242[10] ) );
    nor2_1 \U1652_1_/U2/U5  ( .x(\nchdr_ack[1] ), .a(\net242[9] ), .b(
        \net244[9] ) );
    ao222_2 \U1652_1_/U12/U19/U1/U1  ( .x(\net244[9] ), .a(\net243[9] ), .b(
        csize[1]), .c(\net243[9] ), .d(\net244[9] ), .e(csize[1]), .f(
        \net244[9] ) );
    ao222_2 \U1652_1_/U11/U19/U1/U1  ( .x(\net242[9] ), .a(csize[3]), .b(
        \net243[9] ), .c(csize[3]), .d(\net242[9] ), .e(\net243[9] ), .f(
        \net242[9] ) );
    nor2_1 \U1652_2_/U2/U5  ( .x(\nchdr_ack[2] ), .a(\net242[8] ), .b(
        \net244[8] ) );
    ao222_2 \U1652_2_/U12/U19/U1/U1  ( .x(\net244[8] ), .a(\net243[8] ), .b(
        crnw[0]), .c(\net243[8] ), .d(\net244[8] ), .e(crnw[0]), .f(
        \net244[8] ) );
    ao222_2 \U1652_2_/U11/U19/U1/U1  ( .x(\net242[8] ), .a(crnw[1]), .b(
        \net243[8] ), .c(crnw[1]), .d(\net242[8] ), .e(\net243[8] ), .f(
        \net242[8] ) );
    nor2_1 \U1652_3_/U2/U5  ( .x(\nchdr_ack[3] ), .a(\net242[7] ), .b(
        \net244[7] ) );
    ao222_2 \U1652_3_/U12/U19/U1/U1  ( .x(\net244[7] ), .a(\net243[7] ), .b(
        ctag[0]), .c(\net243[7] ), .d(\net244[7] ), .e(ctag[0]), .f(
        \net244[7] ) );
    ao222_2 \U1652_3_/U11/U19/U1/U1  ( .x(\net242[7] ), .a(ctag[5]), .b(
        \net243[7] ), .c(ctag[5]), .d(\net242[7] ), .e(\net243[7] ), .f(
        \net242[7] ) );
    nor2_1 \U1652_4_/U2/U5  ( .x(\nchdr_ack[4] ), .a(\net242[6] ), .b(
        \net244[6] ) );
    ao222_2 \U1652_4_/U12/U19/U1/U1  ( .x(\net244[6] ), .a(\net243[6] ), .b(
        ctag[1]), .c(\net243[6] ), .d(\net244[6] ), .e(ctag[1]), .f(
        \net244[6] ) );
    ao222_2 \U1652_4_/U11/U19/U1/U1  ( .x(\net242[6] ), .a(ctag[6]), .b(
        \net243[6] ), .c(ctag[6]), .d(\net242[6] ), .e(\net243[6] ), .f(
        \net242[6] ) );
    nor2_1 \U1652_5_/U2/U5  ( .x(\nchdr_ack[5] ), .a(\net242[5] ), .b(
        \net244[5] ) );
    ao222_2 \U1652_5_/U12/U19/U1/U1  ( .x(\net244[5] ), .a(\net243[5] ), .b(
        ctag[2]), .c(\net243[5] ), .d(\net244[5] ), .e(ctag[2]), .f(
        \net244[5] ) );
    ao222_2 \U1652_5_/U11/U19/U1/U1  ( .x(\net242[5] ), .a(ctag[7]), .b(
        \net243[5] ), .c(ctag[7]), .d(\net242[5] ), .e(\net243[5] ), .f(
        \net242[5] ) );
    nor2_1 \U1652_6_/U2/U5  ( .x(\nchdr_ack[6] ), .a(\net242[4] ), .b(
        \net244[4] ) );
    ao222_2 \U1652_6_/U12/U19/U1/U1  ( .x(\net244[4] ), .a(\net243[4] ), .b(
        ctag[3]), .c(\net243[4] ), .d(\net244[4] ), .e(ctag[3]), .f(
        \net244[4] ) );
    ao222_2 \U1652_6_/U11/U19/U1/U1  ( .x(\net242[4] ), .a(ctag[8]), .b(
        \net243[4] ), .c(ctag[8]), .d(\net242[4] ), .e(\net243[4] ), .f(
        \net242[4] ) );
    nor2_1 \U1652_7_/U2/U5  ( .x(\nchdr_ack[7] ), .a(\net242[3] ), .b(
        \net244[3] ) );
    ao222_2 \U1652_7_/U12/U19/U1/U1  ( .x(\net244[3] ), .a(\net243[3] ), .b(
        ctag[4]), .c(\net243[3] ), .d(\net244[3] ), .e(ctag[4]), .f(
        \net244[3] ) );
    ao222_2 \U1652_7_/U11/U19/U1/U1  ( .x(\net242[3] ), .a(ctag[9]), .b(
        \net243[3] ), .c(ctag[9]), .d(\net242[3] ), .e(\net243[3] ), .f(
        \net242[3] ) );
    nor2_1 \U1652_8_/U2/U5  ( .x(\nchdr_ack[8] ), .a(\net242[2] ), .b(
        \net244[2] ) );
    ao222_2 \U1652_8_/U12/U19/U1/U1  ( .x(\net244[2] ), .a(\net243[2] ), .b(
        ccol[0]), .c(\net243[2] ), .d(\net244[2] ), .e(ccol[0]), .f(
        \net244[2] ) );
    ao222_2 \U1652_8_/U11/U19/U1/U1  ( .x(\net242[2] ), .a(ccol[3]), .b(
        \net243[2] ), .c(ccol[3]), .d(\net242[2] ), .e(\net243[2] ), .f(
        \net242[2] ) );
    nor2_1 \U1652_9_/U2/U5  ( .x(\nchdr_ack[9] ), .a(\net242[1] ), .b(
        \net244[1] ) );
    ao222_2 \U1652_9_/U12/U19/U1/U1  ( .x(\net244[1] ), .a(\net243[1] ), .b(
        ccol[1]), .c(\net243[1] ), .d(\net244[1] ), .e(ccol[1]), .f(
        \net244[1] ) );
    ao222_2 \U1652_9_/U11/U19/U1/U1  ( .x(\net242[1] ), .a(ccol[4]), .b(
        \net243[1] ), .c(ccol[4]), .d(\net242[1] ), .e(\net243[1] ), .f(
        \net242[1] ) );
    nor2_1 \U1652_10_/U2/U5  ( .x(\nchdr_ack[10] ), .a(\net242[0] ), .b(
        \net244[0] ) );
    ao222_2 \U1652_10_/U12/U19/U1/U1  ( .x(\net244[0] ), .a(\net243[0] ), .b(
        ccol[2]), .c(\net243[0] ), .d(\net244[0] ), .e(ccol[2]), .f(
        \net244[0] ) );
    ao222_2 \U1652_10_/U11/U19/U1/U1  ( .x(\net242[0] ), .a(ccol[5]), .b(
        \net243[0] ), .c(ccol[5]), .d(\net242[0] ), .e(\net243[0] ), .f(
        \net242[0] ) );
    nor2_1 \U1574_0_/U2/U5  ( .x(\U1574_0_/net231 ), .a(\rhdr_l[5] ), .b(
        \rhdr_h[5] ) );
    and2_1 \U1574_0_/U13/U8  ( .x(\net243[10] ), .a(\U1574_0_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_0_/U12/U19/U1/U1  ( .x(\rhdr_h[5] ), .a(n9), .b(
        \net242[10] ), .c(n9), .d(\rhdr_h[5] ), .e(\net242[10] ), .f(
        \rhdr_h[5] ) );
    ao222_2 \U1574_0_/U11/U19/U1/U1  ( .x(\rhdr_l[5] ), .a(\net244[10] ), .b(
        n8), .c(\net244[10] ), .d(\rhdr_l[5] ), .e(n9), .f(\rhdr_l[5] ) );
    nor2_1 \U1574_1_/U2/U5  ( .x(\U1574_1_/net231 ), .a(\rhdr_l[6] ), .b(
        \rhdr_h[6] ) );
    and2_1 \U1574_1_/U13/U8  ( .x(\net243[9] ), .a(\U1574_1_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_1_/U12/U19/U1/U1  ( .x(\rhdr_h[6] ), .a(n8), .b(\net242[9] 
        ), .c(n7), .d(\rhdr_h[6] ), .e(\net242[9] ), .f(\rhdr_h[6] ) );
    ao222_2 \U1574_1_/U11/U19/U1/U1  ( .x(\rhdr_l[6] ), .a(\net244[9] ), .b(n8
        ), .c(\net244[9] ), .d(\rhdr_l[6] ), .e(n9), .f(\rhdr_l[6] ) );
    nor2_1 \U1574_2_/U2/U5  ( .x(\U1574_2_/net231 ), .a(\rhdr_l[7] ), .b(
        \rhdr_h[7] ) );
    and2_1 \U1574_2_/U13/U8  ( .x(\net243[8] ), .a(\U1574_2_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_2_/U12/U19/U1/U1  ( .x(\rhdr_h[7] ), .a(n7), .b(\net242[8] 
        ), .c(n7), .d(\rhdr_h[7] ), .e(\net242[8] ), .f(\rhdr_h[7] ) );
    ao222_2 \U1574_2_/U11/U19/U1/U1  ( .x(\rhdr_l[7] ), .a(\net244[8] ), .b(n8
        ), .c(\net244[8] ), .d(\rhdr_l[7] ), .e(n9), .f(\rhdr_l[7] ) );
    nor2_1 \U1574_3_/U2/U5  ( .x(\U1574_3_/net231 ), .a(tag_l[0]), .b(tag_h[0]
        ) );
    and2_1 \U1574_3_/U13/U8  ( .x(\net243[7] ), .a(\U1574_3_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_3_/U12/U19/U1/U1  ( .x(tag_h[0]), .a(n9), .b(\net242[7] ), 
        .c(n7), .d(tag_h[0]), .e(\net242[7] ), .f(tag_h[0]) );
    ao222_2 \U1574_3_/U11/U19/U1/U1  ( .x(tag_l[0]), .a(\net244[7] ), .b(n8), 
        .c(\net244[7] ), .d(tag_l[0]), .e(n7), .f(tag_l[0]) );
    nor2_1 \U1574_4_/U2/U5  ( .x(\U1574_4_/net231 ), .a(tag_l[1]), .b(tag_h[1]
        ) );
    and2_1 \U1574_4_/U13/U8  ( .x(\net243[6] ), .a(\U1574_4_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_4_/U12/U19/U1/U1  ( .x(tag_h[1]), .a(n7), .b(\net242[6] ), 
        .c(n7), .d(tag_h[1]), .e(\net242[6] ), .f(tag_h[1]) );
    ao222_2 \U1574_4_/U11/U19/U1/U1  ( .x(tag_l[1]), .a(\net244[6] ), .b(n8), 
        .c(\net244[6] ), .d(tag_l[1]), .e(n7), .f(tag_l[1]) );
    nor2_1 \U1574_5_/U2/U5  ( .x(\U1574_5_/net231 ), .a(tag_l[2]), .b(tag_h[2]
        ) );
    and2_1 \U1574_5_/U13/U8  ( .x(\net243[5] ), .a(\U1574_5_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_5_/U12/U19/U1/U1  ( .x(tag_h[2]), .a(n8), .b(\net242[5] ), 
        .c(n7), .d(tag_h[2]), .e(\net242[5] ), .f(tag_h[2]) );
    ao222_2 \U1574_5_/U11/U19/U1/U1  ( .x(tag_l[2]), .a(\net244[5] ), .b(n8), 
        .c(\net244[5] ), .d(tag_l[2]), .e(n9), .f(tag_l[2]) );
    nor2_1 \U1574_6_/U2/U5  ( .x(\U1574_6_/net231 ), .a(tag_l[3]), .b(tag_h[3]
        ) );
    and2_1 \U1574_6_/U13/U8  ( .x(\net243[4] ), .a(\U1574_6_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_6_/U12/U19/U1/U1  ( .x(tag_h[3]), .a(n7), .b(\net242[4] ), 
        .c(n9), .d(tag_h[3]), .e(\net242[4] ), .f(tag_h[3]) );
    ao222_2 \U1574_6_/U11/U19/U1/U1  ( .x(tag_l[3]), .a(\net244[4] ), .b(n8), 
        .c(\net244[4] ), .d(tag_l[3]), .e(n7), .f(tag_l[3]) );
    nor2_1 \U1574_7_/U2/U5  ( .x(\U1574_7_/net231 ), .a(tag_l[4]), .b(tag_h[4]
        ) );
    and2_1 \U1574_7_/U13/U8  ( .x(\net243[3] ), .a(\U1574_7_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_7_/U12/U19/U1/U1  ( .x(tag_h[4]), .a(n7), .b(\net242[3] ), 
        .c(n9), .d(tag_h[4]), .e(\net242[3] ), .f(tag_h[4]) );
    ao222_2 \U1574_7_/U11/U19/U1/U1  ( .x(tag_l[4]), .a(\net244[3] ), .b(n8), 
        .c(\net244[3] ), .d(tag_l[4]), .e(n7), .f(tag_l[4]) );
    nor2_1 \U1574_8_/U2/U5  ( .x(\U1574_8_/net231 ), .a(\rhdr_l[13] ), .b(
        \rhdr_h[13] ) );
    and2_1 \U1574_8_/U13/U8  ( .x(\net243[2] ), .a(\U1574_8_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_8_/U12/U19/U1/U1  ( .x(\rhdr_h[13] ), .a(n8), .b(
        \net242[2] ), .c(n9), .d(\rhdr_h[13] ), .e(\net242[2] ), .f(
        \rhdr_h[13] ) );
    ao222_2 \U1574_8_/U11/U19/U1/U1  ( .x(\rhdr_l[13] ), .a(\net244[2] ), .b(
        n8), .c(\net244[2] ), .d(\rhdr_l[13] ), .e(n7), .f(\rhdr_l[13] ) );
    nor2_1 \U1574_9_/U2/U5  ( .x(\U1574_9_/net231 ), .a(\rhdr_l[14] ), .b(
        \rhdr_h[14] ) );
    and2_1 \U1574_9_/U13/U8  ( .x(\net243[1] ), .a(\U1574_9_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_9_/U12/U19/U1/U1  ( .x(\rhdr_h[14] ), .a(n9), .b(
        \net242[1] ), .c(n7), .d(\rhdr_h[14] ), .e(\net242[1] ), .f(
        \rhdr_h[14] ) );
    ao222_2 \U1574_9_/U11/U19/U1/U1  ( .x(\rhdr_l[14] ), .a(\net244[1] ), .b(
        n8), .c(\net244[1] ), .d(\rhdr_l[14] ), .e(n9), .f(\rhdr_l[14] ) );
    nor2_1 \U1574_10_/U2/U5  ( .x(\U1574_10_/net231 ), .a(\rhdr_l[15] ), .b(
        \rhdr_h[15] ) );
    and2_1 \U1574_10_/U13/U8  ( .x(\net243[0] ), .a(\U1574_10_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_10_/U12/U19/U1/U1  ( .x(\rhdr_h[15] ), .a(n9), .b(
        \net242[0] ), .c(n9), .d(\rhdr_h[15] ), .e(\net242[0] ), .f(
        \rhdr_h[15] ) );
    ao222_2 \U1574_10_/U11/U19/U1/U1  ( .x(\rhdr_l[15] ), .a(\net244[0] ), .b(
        n8), .c(\net244[0] ), .d(\rhdr_l[15] ), .e(n9), .f(\rhdr_l[15] ) );
    buf_1 U1 ( .x(csize[0]), .a(n14) );
    buf_1 U2 ( .x(csize[1]), .a(n13) );
    buf_1 U3 ( .x(csize[3]), .a(n12) );
    buf_1 U4 ( .x(crnw[0]), .a(n11) );
    buf_1 U5 ( .x(crnw[1]), .a(n10) );
    inv_5 U6 ( .x(n6), .a(net265) );
    buf_3 U7 ( .x(nbreset), .a(nReset) );
    buf_3 U8 ( .x(n7), .a(net248) );
    buf_3 U9 ( .x(n9), .a(net248) );
    buf_3 U10 ( .x(n8), .a(net248) );
    nor2_1 U11 ( .x(net248), .a(net265), .b(rhdrack) );
endmodule


module chain_selement_ga_19 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_18 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[1] , \c[0] ;
    chain_selement_ga_19 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_20 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_19 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[1] , \c[0] ;
    chain_selement_ga_20 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_21 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_20 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[1] , \c[0] , n1, n2;
    chain_selement_ga_21 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        n2), .e(n2) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(n2), .b(r[0]), .c(n2), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(n2), .b(r[1]), .c(n2), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
    inv_0 U1 ( .x(n1), .a(e[0]) );
    inv_2 U2 ( .x(n2), .a(n1) );
endmodule


module chain_selement_ga_76 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module resp_route_tx_dmem ( o, rtxack, e_h, e_l, noa, r_h, r_l, rtxreq );
output [4:0] o;
input  [2:0] e_h;
input  [2:0] e_l;
input  [2:0] r_h;
input  [2:0] r_l;
input  noa, rtxreq;
output rtxack;
    wire \r2[2] , \r2[1] , \r2[0] , \r1[2] , \r1[1] , \r1[0] , \r0[2] , 
        \r0[1] , \r0[0] , \last[0] , \last[1] , \last[2] , \last[3] , 
        \net72[0] , \net72[1] , net56, net106, net103, eopsym, net87, net66, 
        net84, net77, \I8/nb , \I8/na , \I11/n5 , \I11/n1 , \I11/n2 , \I11/n3 , 
        \I11/n4 , \I7_0_/U25/U1/clr , \I7_0_/U25/U1/ob , \I7_1_/U25/U1/clr , 
        \I7_1_/U25/U1/ob ;
    assign o[3] = 1'b0;
    assign o[2] = 1'b0;
    chain_selement_ga_76 I9 ( .Aa(\last[0] ), .Br(eopsym), .Ar(net87), .Ba(
        net66) );
    route_symbol_19 I2 ( .o({\r1[2] , \r1[1] , \r1[0] }), .txack(net84), 
        .txack_last(\last[2] ), .e({e_h[1], e_l[1]}), .oa(net66), .r({r_h[1], 
        r_l[1]}), .txreq(net77) );
    route_symbol_20 I3 ( .o({\r0[2] , \r0[1] , \r0[0] }), .txack(net87), 
        .txack_last(\last[1] ), .e({e_h[0], e_l[0]}), .oa(net66), .r({r_h[0], 
        r_l[0]}), .txreq(net84) );
    route_symbol_18 I1 ( .o({\r2[2] , \r2[1] , \r2[0] }), .txack(net77), 
        .txack_last(\last[3] ), .e({e_h[2], e_l[2]}), .oa(net66), .r({r_h[2], 
        r_l[2]}), .txreq(rtxreq) );
    nor2_1 \I5/U5  ( .x(net106), .a(eopsym), .b(\r2[2] ) );
    nor2_1 \I16/U5  ( .x(net103), .a(\r1[2] ), .b(\r0[2] ) );
    or2_1 \I14_0_/U12  ( .x(\net72[1] ), .a(\r2[0] ), .b(\r1[0] ) );
    or2_1 \I14_1_/U12  ( .x(\net72[0] ), .a(\r2[1] ), .b(\r1[1] ) );
    nor3_1 \I8/U27  ( .x(\I8/nb ), .a(o[4]), .b(o[3]), .c(o[2]) );
    nor2_1 \I8/U26  ( .x(\I8/na ), .a(o[1]), .b(o[0]) );
    nand2_2 \I8/U29  ( .x(net66), .a(\I8/nb ), .b(\I8/na ) );
    and4_1 \I11/U16  ( .x(\I11/n5 ), .a(\I11/n1 ), .b(\I11/n2 ), .c(\I11/n3 ), 
        .d(\I11/n4 ) );
    inv_1 \I11/U1  ( .x(\I11/n1 ), .a(\last[3] ) );
    inv_1 \I11/U2  ( .x(\I11/n2 ), .a(\last[2] ) );
    inv_1 \I11/U3  ( .x(\I11/n3 ), .a(\last[1] ) );
    inv_1 \I11/U4  ( .x(\I11/n4 ), .a(\last[0] ) );
    inv_1 \I11/U5  ( .x(rtxack), .a(\I11/n5 ) );
    nand2_1 \I17/U5  ( .x(net56), .a(net106), .b(net103) );
    ao222_1 \I15/U18/U1/U1  ( .x(o[4]), .a(noa), .b(net56), .c(noa), .d(o[4]), 
        .e(net56), .f(o[4]) );
    oa31_1 \I7_0_/U25/U1/Uclr  ( .x(\I7_0_/U25/U1/clr ), .a(noa), .b(\r0[0] ), 
        .c(\net72[1] ), .d(o[0]) );
    oaoi211_1 \I7_0_/U25/U1/Uaoi  ( .x(\I7_0_/U25/U1/ob ), .a(\r0[0] ), .b(
        \net72[1] ), .c(noa), .d(\I7_0_/U25/U1/clr ) );
    inv_2 \I7_0_/U25/U1/Ui  ( .x(o[0]), .a(\I7_0_/U25/U1/ob ) );
    oa31_1 \I7_1_/U25/U1/Uclr  ( .x(\I7_1_/U25/U1/clr ), .a(noa), .b(\r0[1] ), 
        .c(\net72[0] ), .d(o[1]) );
    oaoi211_1 \I7_1_/U25/U1/Uaoi  ( .x(\I7_1_/U25/U1/ob ), .a(\r0[1] ), .b(
        \net72[0] ), .c(noa), .d(\I7_1_/U25/U1/clr ) );
    inv_2 \I7_1_/U25/U1/Ui  ( .x(o[1]), .a(\I7_1_/U25/U1/ob ) );
endmodule


module matched_delay_cp2slave_resp_dmem ( x, a );
input  a;
output x;
    buf_1 I1 ( .x(x), .a(a) );
endmodule


module matched_delay_cp2slave_comdmem ( x, a );
input  a;
output x;
    buf_1 I1 ( .x(x), .a(a) );
endmodule


module sr2dr_word_8 ( i, req, h, l );
input  [31:0] i;
output [31:0] h;
output [31:0] l;
input  req;
    wire \U31/nl , \U31/ni , \U31/nh , \U30/nl , \U30/ni , \U30/nh , \U29/nl , 
        \U29/ni , \U29/nh , \U28/nl , \U28/ni , \U28/nh , \U27/nl , \U27/ni , 
        \U27/nh , \U26/nl , \U26/ni , \U26/nh , \U25/nl , \U25/ni , \U25/nh , 
        \U24/nl , \U24/ni , \U24/nh , \U23/nl , \U23/ni , \U23/nh , \U22/nl , 
        \U22/ni , \U22/nh , \U21/nl , \U21/ni , \U21/nh , \U20/nl , \U20/ni , 
        \U20/nh , \U19/nl , \U19/ni , \U19/nh , \U18/nl , \U18/ni , \U18/nh , 
        \U17/nl , \U17/ni , \U17/nh , \U16/nl , \U16/ni , \U16/nh , \U15/nl , 
        \U15/ni , \U15/nh , \U14/nl , \U14/ni , \U14/nh , \U13/nl , \U13/ni , 
        \U13/nh , \U12/nl , \U12/ni , \U12/nh , \U11/nl , \U11/ni , \U11/nh , 
        \U10/nl , \U10/ni , \U10/nh , \U9/nl , \U9/ni , \U9/nh , \U8/nl , 
        \U8/ni , \U8/nh , \U7/nl , \U7/ni , \U7/nh , \U6/nl , \U6/ni , \U6/nh , 
        \U5/nl , \U5/ni , \U5/nh , \U4/nl , \U4/ni , \U4/nh , \U3/nl , \U3/ni , 
        \U3/nh , \U2/nl , \U2/ni , \U2/nh , \U1/nl , \U1/ni , \U1/nh , \U0/nl , 
        \U0/ni , \U0/nh , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
    inv_1 \U31/Uii  ( .x(\U31/ni ), .a(i[31]) );
    inv_1 \U31/Uih  ( .x(\U31/nh ), .a(h[31]) );
    inv_1 \U31/Uil  ( .x(\U31/nl ), .a(l[31]) );
    ao23_1 \U31/Ucl/U1/U1  ( .x(l[31]), .a(n9), .b(l[31]), .c(n1), .d(\U31/ni 
        ), .e(\U31/nh ) );
    ao23_1 \U31/Uch/U1/U1  ( .x(h[31]), .a(n9), .b(h[31]), .c(n2), .d(i[31]), 
        .e(\U31/nl ) );
    inv_1 \U30/Uii  ( .x(\U30/ni ), .a(i[30]) );
    inv_1 \U30/Uih  ( .x(\U30/nh ), .a(h[30]) );
    inv_1 \U30/Uil  ( .x(\U30/nl ), .a(l[30]) );
    ao23_1 \U30/Ucl/U1/U1  ( .x(l[30]), .a(n8), .b(l[30]), .c(n1), .d(\U30/ni 
        ), .e(\U30/nh ) );
    ao23_1 \U30/Uch/U1/U1  ( .x(h[30]), .a(n8), .b(h[30]), .c(n1), .d(i[30]), 
        .e(\U30/nl ) );
    inv_1 \U29/Uii  ( .x(\U29/ni ), .a(i[29]) );
    inv_1 \U29/Uih  ( .x(\U29/nh ), .a(h[29]) );
    inv_1 \U29/Uil  ( .x(\U29/nl ), .a(l[29]) );
    ao23_1 \U29/Ucl/U1/U1  ( .x(l[29]), .a(n8), .b(l[29]), .c(n1), .d(\U29/ni 
        ), .e(\U29/nh ) );
    ao23_1 \U29/Uch/U1/U1  ( .x(h[29]), .a(n8), .b(h[29]), .c(n2), .d(i[29]), 
        .e(\U29/nl ) );
    inv_1 \U28/Uii  ( .x(\U28/ni ), .a(i[28]) );
    inv_1 \U28/Uih  ( .x(\U28/nh ), .a(h[28]) );
    inv_1 \U28/Uil  ( .x(\U28/nl ), .a(l[28]) );
    ao23_1 \U28/Ucl/U1/U1  ( .x(l[28]), .a(n8), .b(l[28]), .c(n2), .d(\U28/ni 
        ), .e(\U28/nh ) );
    ao23_1 \U28/Uch/U1/U1  ( .x(h[28]), .a(n8), .b(h[28]), .c(n2), .d(i[28]), 
        .e(\U28/nl ) );
    inv_1 \U27/Uii  ( .x(\U27/ni ), .a(i[27]) );
    inv_1 \U27/Uih  ( .x(\U27/nh ), .a(h[27]) );
    inv_1 \U27/Uil  ( .x(\U27/nl ), .a(l[27]) );
    ao23_1 \U27/Ucl/U1/U1  ( .x(l[27]), .a(n8), .b(l[27]), .c(n2), .d(\U27/ni 
        ), .e(\U27/nh ) );
    ao23_1 \U27/Uch/U1/U1  ( .x(h[27]), .a(n8), .b(h[27]), .c(n2), .d(i[27]), 
        .e(\U27/nl ) );
    inv_1 \U26/Uii  ( .x(\U26/ni ), .a(i[26]) );
    inv_1 \U26/Uih  ( .x(\U26/nh ), .a(h[26]) );
    inv_1 \U26/Uil  ( .x(\U26/nl ), .a(l[26]) );
    ao23_1 \U26/Ucl/U1/U1  ( .x(l[26]), .a(n7), .b(l[26]), .c(n2), .d(\U26/ni 
        ), .e(\U26/nh ) );
    ao23_1 \U26/Uch/U1/U1  ( .x(h[26]), .a(n7), .b(h[26]), .c(n4), .d(i[26]), 
        .e(\U26/nl ) );
    inv_1 \U25/Uii  ( .x(\U25/ni ), .a(i[25]) );
    inv_1 \U25/Uih  ( .x(\U25/nh ), .a(h[25]) );
    inv_1 \U25/Uil  ( .x(\U25/nl ), .a(l[25]) );
    ao23_1 \U25/Ucl/U1/U1  ( .x(l[25]), .a(n7), .b(l[25]), .c(n4), .d(\U25/ni 
        ), .e(\U25/nh ) );
    ao23_1 \U25/Uch/U1/U1  ( .x(h[25]), .a(n7), .b(h[25]), .c(n4), .d(i[25]), 
        .e(\U25/nl ) );
    inv_1 \U24/Uii  ( .x(\U24/ni ), .a(i[24]) );
    inv_1 \U24/Uih  ( .x(\U24/nh ), .a(h[24]) );
    inv_1 \U24/Uil  ( .x(\U24/nl ), .a(l[24]) );
    ao23_1 \U24/Ucl/U1/U1  ( .x(l[24]), .a(n7), .b(l[24]), .c(n4), .d(\U24/ni 
        ), .e(\U24/nh ) );
    ao23_1 \U24/Uch/U1/U1  ( .x(h[24]), .a(n7), .b(h[24]), .c(n4), .d(i[24]), 
        .e(\U24/nl ) );
    inv_1 \U23/Uii  ( .x(\U23/ni ), .a(i[23]) );
    inv_1 \U23/Uih  ( .x(\U23/nh ), .a(h[23]) );
    inv_1 \U23/Uil  ( .x(\U23/nl ), .a(l[23]) );
    ao23_1 \U23/Ucl/U1/U1  ( .x(l[23]), .a(n7), .b(l[23]), .c(n3), .d(\U23/ni 
        ), .e(\U23/nh ) );
    ao23_1 \U23/Uch/U1/U1  ( .x(h[23]), .a(n7), .b(h[23]), .c(n3), .d(i[23]), 
        .e(\U23/nl ) );
    inv_1 \U22/Uii  ( .x(\U22/ni ), .a(i[22]) );
    inv_1 \U22/Uih  ( .x(\U22/nh ), .a(h[22]) );
    inv_1 \U22/Uil  ( .x(\U22/nl ), .a(l[22]) );
    ao23_1 \U22/Ucl/U1/U1  ( .x(l[22]), .a(n6), .b(l[22]), .c(n3), .d(\U22/ni 
        ), .e(\U22/nh ) );
    ao23_1 \U22/Uch/U1/U1  ( .x(h[22]), .a(n6), .b(h[22]), .c(n3), .d(i[22]), 
        .e(\U22/nl ) );
    inv_1 \U21/Uii  ( .x(\U21/ni ), .a(i[21]) );
    inv_1 \U21/Uih  ( .x(\U21/nh ), .a(h[21]) );
    inv_1 \U21/Uil  ( .x(\U21/nl ), .a(l[21]) );
    ao23_1 \U21/Ucl/U1/U1  ( .x(l[21]), .a(n6), .b(l[21]), .c(n3), .d(\U21/ni 
        ), .e(\U21/nh ) );
    ao23_1 \U21/Uch/U1/U1  ( .x(h[21]), .a(n6), .b(h[21]), .c(n3), .d(i[21]), 
        .e(\U21/nl ) );
    inv_1 \U20/Uii  ( .x(\U20/ni ), .a(i[20]) );
    inv_1 \U20/Uih  ( .x(\U20/nh ), .a(h[20]) );
    inv_1 \U20/Uil  ( .x(\U20/nl ), .a(l[20]) );
    ao23_1 \U20/Ucl/U1/U1  ( .x(l[20]), .a(n6), .b(l[20]), .c(n5), .d(\U20/ni 
        ), .e(\U20/nh ) );
    ao23_1 \U20/Uch/U1/U1  ( .x(h[20]), .a(n6), .b(h[20]), .c(n4), .d(i[20]), 
        .e(\U20/nl ) );
    inv_1 \U19/Uii  ( .x(\U19/ni ), .a(i[19]) );
    inv_1 \U19/Uih  ( .x(\U19/nh ), .a(h[19]) );
    inv_1 \U19/Uil  ( .x(\U19/nl ), .a(l[19]) );
    ao23_1 \U19/Ucl/U1/U1  ( .x(l[19]), .a(n6), .b(l[19]), .c(n4), .d(\U19/ni 
        ), .e(\U19/nh ) );
    ao23_1 \U19/Uch/U1/U1  ( .x(h[19]), .a(n6), .b(h[19]), .c(n4), .d(i[19]), 
        .e(\U19/nl ) );
    inv_1 \U18/Uii  ( .x(\U18/ni ), .a(i[18]) );
    inv_1 \U18/Uih  ( .x(\U18/nh ), .a(h[18]) );
    inv_1 \U18/Uil  ( .x(\U18/nl ), .a(l[18]) );
    ao23_1 \U18/Ucl/U1/U1  ( .x(l[18]), .a(n5), .b(l[18]), .c(n5), .d(\U18/ni 
        ), .e(\U18/nh ) );
    ao23_1 \U18/Uch/U1/U1  ( .x(h[18]), .a(n5), .b(h[18]), .c(n5), .d(i[18]), 
        .e(\U18/nl ) );
    inv_1 \U17/Uii  ( .x(\U17/ni ), .a(i[17]) );
    inv_1 \U17/Uih  ( .x(\U17/nh ), .a(h[17]) );
    inv_1 \U17/Uil  ( .x(\U17/nl ), .a(l[17]) );
    ao23_1 \U17/Ucl/U1/U1  ( .x(l[17]), .a(n6), .b(l[17]), .c(n5), .d(\U17/ni 
        ), .e(\U17/nh ) );
    ao23_1 \U17/Uch/U1/U1  ( .x(h[17]), .a(n7), .b(h[17]), .c(n4), .d(i[17]), 
        .e(\U17/nl ) );
    inv_1 \U16/Uii  ( .x(\U16/ni ), .a(i[16]) );
    inv_1 \U16/Uih  ( .x(\U16/nh ), .a(h[16]) );
    inv_1 \U16/Uil  ( .x(\U16/nl ), .a(l[16]) );
    ao23_1 \U16/Ucl/U1/U1  ( .x(l[16]), .a(n9), .b(l[16]), .c(n3), .d(\U16/ni 
        ), .e(\U16/nh ) );
    ao23_1 \U16/Uch/U1/U1  ( .x(h[16]), .a(n9), .b(h[16]), .c(n1), .d(i[16]), 
        .e(\U16/nl ) );
    inv_1 \U15/Uii  ( .x(\U15/ni ), .a(i[15]) );
    inv_1 \U15/Uih  ( .x(\U15/nh ), .a(h[15]) );
    inv_1 \U15/Uil  ( .x(\U15/nl ), .a(l[15]) );
    ao23_1 \U15/Ucl/U1/U1  ( .x(l[15]), .a(n8), .b(l[15]), .c(n1), .d(\U15/ni 
        ), .e(\U15/nh ) );
    ao23_1 \U15/Uch/U1/U1  ( .x(h[15]), .a(n7), .b(h[15]), .c(n1), .d(i[15]), 
        .e(\U15/nl ) );
    inv_1 \U14/Uii  ( .x(\U14/ni ), .a(i[14]) );
    inv_1 \U14/Uih  ( .x(\U14/nh ), .a(h[14]) );
    inv_1 \U14/Uil  ( .x(\U14/nl ), .a(l[14]) );
    ao23_1 \U14/Ucl/U1/U1  ( .x(l[14]), .a(n6), .b(l[14]), .c(n1), .d(\U14/ni 
        ), .e(\U14/nh ) );
    ao23_1 \U14/Uch/U1/U1  ( .x(h[14]), .a(n6), .b(h[14]), .c(n3), .d(i[14]), 
        .e(\U14/nl ) );
    inv_1 \U13/Uii  ( .x(\U13/ni ), .a(i[13]) );
    inv_1 \U13/Uih  ( .x(\U13/nh ), .a(h[13]) );
    inv_1 \U13/Uil  ( .x(\U13/nl ), .a(l[13]) );
    ao23_1 \U13/Ucl/U1/U1  ( .x(l[13]), .a(n6), .b(l[13]), .c(n4), .d(\U13/ni 
        ), .e(\U13/nh ) );
    ao23_1 \U13/Uch/U1/U1  ( .x(h[13]), .a(n6), .b(h[13]), .c(n4), .d(i[13]), 
        .e(\U13/nl ) );
    inv_1 \U12/Uii  ( .x(\U12/ni ), .a(i[12]) );
    inv_1 \U12/Uih  ( .x(\U12/nh ), .a(h[12]) );
    inv_1 \U12/Uil  ( .x(\U12/nl ), .a(l[12]) );
    ao23_1 \U12/Ucl/U1/U1  ( .x(l[12]), .a(n5), .b(l[12]), .c(n4), .d(\U12/ni 
        ), .e(\U12/nh ) );
    ao23_1 \U12/Uch/U1/U1  ( .x(h[12]), .a(n5), .b(h[12]), .c(n4), .d(i[12]), 
        .e(\U12/nl ) );
    inv_1 \U11/Uii  ( .x(\U11/ni ), .a(i[11]) );
    inv_1 \U11/Uih  ( .x(\U11/nh ), .a(h[11]) );
    inv_1 \U11/Uil  ( .x(\U11/nl ), .a(l[11]) );
    ao23_1 \U11/Ucl/U1/U1  ( .x(l[11]), .a(n5), .b(l[11]), .c(n4), .d(\U11/ni 
        ), .e(\U11/nh ) );
    ao23_1 \U11/Uch/U1/U1  ( .x(h[11]), .a(n5), .b(h[11]), .c(n4), .d(i[11]), 
        .e(\U11/nl ) );
    inv_1 \U10/Uii  ( .x(\U10/ni ), .a(i[10]) );
    inv_1 \U10/Uih  ( .x(\U10/nh ), .a(h[10]) );
    inv_1 \U10/Uil  ( .x(\U10/nl ), .a(l[10]) );
    ao23_1 \U10/Ucl/U1/U1  ( .x(l[10]), .a(n5), .b(l[10]), .c(n3), .d(\U10/ni 
        ), .e(\U10/nh ) );
    ao23_1 \U10/Uch/U1/U1  ( .x(h[10]), .a(n5), .b(h[10]), .c(n3), .d(i[10]), 
        .e(\U10/nl ) );
    inv_1 \U9/Uii  ( .x(\U9/ni ), .a(i[9]) );
    inv_1 \U9/Uih  ( .x(\U9/nh ), .a(h[9]) );
    inv_1 \U9/Uil  ( .x(\U9/nl ), .a(l[9]) );
    ao23_1 \U9/Ucl/U1/U1  ( .x(l[9]), .a(n5), .b(l[9]), .c(n3), .d(\U9/ni ), 
        .e(\U9/nh ) );
    ao23_1 \U9/Uch/U1/U1  ( .x(h[9]), .a(n5), .b(h[9]), .c(n3), .d(i[9]), .e(
        \U9/nl ) );
    inv_1 \U8/Uii  ( .x(\U8/ni ), .a(i[8]) );
    inv_1 \U8/Uih  ( .x(\U8/nh ), .a(h[8]) );
    inv_1 \U8/Uil  ( .x(\U8/nl ), .a(l[8]) );
    ao23_1 \U8/Ucl/U1/U1  ( .x(l[8]), .a(n5), .b(l[8]), .c(n3), .d(\U8/ni ), 
        .e(\U8/nh ) );
    ao23_1 \U8/Uch/U1/U1  ( .x(h[8]), .a(n5), .b(h[8]), .c(n3), .d(i[8]), .e(
        \U8/nl ) );
    inv_1 \U7/Uii  ( .x(\U7/ni ), .a(i[7]) );
    inv_1 \U7/Uih  ( .x(\U7/nh ), .a(h[7]) );
    inv_1 \U7/Uil  ( .x(\U7/nl ), .a(l[7]) );
    ao23_1 \U7/Ucl/U1/U1  ( .x(l[7]), .a(n7), .b(l[7]), .c(n3), .d(\U7/ni ), 
        .e(\U7/nh ) );
    ao23_1 \U7/Uch/U1/U1  ( .x(h[7]), .a(n7), .b(h[7]), .c(n2), .d(i[7]), .e(
        \U7/nl ) );
    inv_1 \U6/Uii  ( .x(\U6/ni ), .a(i[6]) );
    inv_1 \U6/Uih  ( .x(\U6/nh ), .a(h[6]) );
    inv_1 \U6/Uil  ( .x(\U6/nl ), .a(l[6]) );
    ao23_1 \U6/Ucl/U1/U1  ( .x(l[6]), .a(n7), .b(l[6]), .c(n2), .d(\U6/ni ), 
        .e(\U6/nh ) );
    ao23_1 \U6/Uch/U1/U1  ( .x(h[6]), .a(n7), .b(h[6]), .c(n2), .d(i[6]), .e(
        \U6/nl ) );
    inv_1 \U5/Uii  ( .x(\U5/ni ), .a(i[5]) );
    inv_1 \U5/Uih  ( .x(\U5/nh ), .a(h[5]) );
    inv_1 \U5/Uil  ( .x(\U5/nl ), .a(l[5]) );
    ao23_1 \U5/Ucl/U1/U1  ( .x(l[5]), .a(n7), .b(l[5]), .c(n2), .d(\U5/ni ), 
        .e(\U5/nh ) );
    ao23_1 \U5/Uch/U1/U1  ( .x(h[5]), .a(n7), .b(h[5]), .c(n2), .d(i[5]), .e(
        \U5/nl ) );
    inv_1 \U4/Uii  ( .x(\U4/ni ), .a(i[4]) );
    inv_1 \U4/Uih  ( .x(\U4/nh ), .a(h[4]) );
    inv_1 \U4/Uil  ( .x(\U4/nl ), .a(l[4]) );
    ao23_1 \U4/Ucl/U1/U1  ( .x(l[4]), .a(n6), .b(l[4]), .c(n2), .d(\U4/ni ), 
        .e(\U4/nh ) );
    ao23_1 \U4/Uch/U1/U1  ( .x(h[4]), .a(n6), .b(h[4]), .c(n2), .d(i[4]), .e(
        \U4/nl ) );
    inv_1 \U3/Uii  ( .x(\U3/ni ), .a(i[3]) );
    inv_1 \U3/Uih  ( .x(\U3/nh ), .a(h[3]) );
    inv_1 \U3/Uil  ( .x(\U3/nl ), .a(l[3]) );
    ao23_1 \U3/Ucl/U1/U1  ( .x(l[3]), .a(n6), .b(l[3]), .c(n2), .d(\U3/ni ), 
        .e(\U3/nh ) );
    ao23_1 \U3/Uch/U1/U1  ( .x(h[3]), .a(n8), .b(h[3]), .c(n1), .d(i[3]), .e(
        \U3/nl ) );
    inv_1 \U2/Uii  ( .x(\U2/ni ), .a(i[2]) );
    inv_1 \U2/Uih  ( .x(\U2/nh ), .a(h[2]) );
    inv_1 \U2/Uil  ( .x(\U2/nl ), .a(l[2]) );
    ao23_1 \U2/Ucl/U1/U1  ( .x(l[2]), .a(n8), .b(l[2]), .c(n1), .d(\U2/ni ), 
        .e(\U2/nh ) );
    ao23_1 \U2/Uch/U1/U1  ( .x(h[2]), .a(n8), .b(h[2]), .c(n1), .d(i[2]), .e(
        \U2/nl ) );
    inv_1 \U1/Uii  ( .x(\U1/ni ), .a(i[1]) );
    inv_1 \U1/Uih  ( .x(\U1/nh ), .a(h[1]) );
    inv_1 \U1/Uil  ( .x(\U1/nl ), .a(l[1]) );
    ao23_1 \U1/Ucl/U1/U1  ( .x(l[1]), .a(n8), .b(l[1]), .c(n1), .d(\U1/ni ), 
        .e(\U1/nh ) );
    ao23_1 \U1/Uch/U1/U1  ( .x(h[1]), .a(n8), .b(h[1]), .c(n1), .d(i[1]), .e(
        \U1/nl ) );
    inv_1 \U0/Uii  ( .x(\U0/ni ), .a(i[0]) );
    inv_1 \U0/Uih  ( .x(\U0/nh ), .a(h[0]) );
    inv_1 \U0/Uil  ( .x(\U0/nl ), .a(l[0]) );
    ao23_1 \U0/Ucl/U1/U1  ( .x(l[0]), .a(n8), .b(l[0]), .c(n1), .d(\U0/ni ), 
        .e(\U0/nh ) );
    ao23_1 \U0/Uch/U1/U1  ( .x(h[0]), .a(n8), .b(h[0]), .c(n1), .d(i[0]), .e(
        \U0/nl ) );
    buf_16 U1 ( .x(n1), .a(n12) );
    buf_16 U2 ( .x(n2), .a(n12) );
    buf_16 U3 ( .x(n3), .a(n12) );
    buf_16 U4 ( .x(n4), .a(n11) );
    buf_16 U5 ( .x(n5), .a(n11) );
    buf_16 U6 ( .x(n6), .a(n11) );
    buf_16 U7 ( .x(n7), .a(n10) );
    buf_16 U8 ( .x(n8), .a(n10) );
    buf_16 U9 ( .x(n9), .a(n10) );
    buf_16 U10 ( .x(n10), .a(req) );
    buf_16 U11 ( .x(n11), .a(req) );
    buf_16 U12 ( .x(n12), .a(req) );
endmodule


module cp2slave_dmem ( tc_seq, tc_size, tc_itag, tc_wd, tc_lock, tc_a, tc_rnw, 
    tc_ok, tc_defer, tc_slow, tc_ack, req_in, ts_i, st_i, we_i, mult_i, adr_i, 
    dat_i, seq_i, prd_i, sel_i, ack_in, tr_rd, tr_err, tr_size, tr_ack, tr_rnw, 
    req_out, dat_o, err_o, rty_o, acc_o, sel_o, mult_o, rt_o, ack_out, reset
     );
input  [1:0] tc_seq;
input  [3:0] tc_size;
input  [9:0] tc_itag;
input  [63:0] tc_wd;
input  [1:0] tc_lock;
input  [63:0] tc_a;
input  [1:0] tc_rnw;
output [2:0] ts_i;
output [4:0] st_i;
output [31:0] adr_i;
output [31:0] dat_i;
output [3:0] sel_i;
output [63:0] tr_rd;
output [1:0] tr_err;
output [3:0] tr_size;
output [1:0] tr_rnw;
input  [31:0] dat_o;
input  [3:0] sel_o;
input  [4:0] rt_o;
input  ack_in, tr_ack, req_out, err_o, rty_o, acc_o, mult_o, reset;
output tc_ok, tc_defer, tc_slow, tc_ack, req_in, we_i, mult_i, seq_i, prd_i, 
    ack_out;
    wire \tc_a[60] , \tc_a[58] , \tc_wd[63] , \tc_wd[62] , \tc_wd[61] , 
        \tc_wd[60] , \tc_wd[59] , \tc_wd[58] , \tc_wd[56] , \tc_wd[55] , 
        \tc_wd[54] , \tc_wd[53] , \tc_wd[52] , \tc_wd[51] , \tc_wd[50] , 
        \tc_wd[49] , \tc_wd[48] , \tc_wd[47] , \tc_wd[46] , \tc_wd[45] , 
        \tc_wd[44] , \tc_wd[43] , \tc_wd[40] , \tc_wd[39] , \tc_wd[38] , 
        \tc_wd[36] , \tc_wd[32] , \sel_i[2] , n121, n122, n123, n124, n125, 
        n126, n127, n128, n129, n130, n135, n136, n137, n141, n142, n180, n181, 
        n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, 
        n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, 
        n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, 
        n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
        n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, 
        n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, 
        n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, 
        n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, 
        n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, 
        n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, 
        n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, 
        n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, 
        n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, 
        n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, 
        n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, 
        n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, 
        n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, 
        n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, 
        n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
        n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
        n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
        n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
        n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
        n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
        n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
        n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
        n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
        n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
        n518, n519, n520, n521, n522, n523, n524, n525, n529, n530, n531, n532, 
        n3, n4, n5, complb1, complb0, comp_basic, complw1, complw0, comp_wd, 
        all_w, all_r, respond, _24_net_, _25_net_, _26_net_, req_out_delayed, 
        req_in_i, \cg_all_w/__tmp99/loop , \Usze1/nl , \Usze1/ni , \Usze1/nh , 
        \Usze0/nl , \Usze0/ni , \Usze0/nh , \Urnw/nl , \Urnw/ni , \Urnw/nh , 
        \Uerr/nl , \Uerr/ni , \Uerr/nh , n1, n2;
    assign \tc_wd[63]  = tc_wd[63];
    assign \tc_wd[62]  = tc_wd[62];
    assign \tc_wd[61]  = tc_wd[61];
    assign \tc_wd[60]  = tc_wd[60];
    assign \tc_wd[59]  = tc_wd[59];
    assign \tc_wd[58]  = tc_wd[58];
    assign \tc_wd[56]  = tc_wd[56];
    assign \tc_wd[55]  = tc_wd[55];
    assign \tc_wd[54]  = tc_wd[54];
    assign \tc_wd[53]  = tc_wd[53];
    assign \tc_wd[52]  = tc_wd[52];
    assign \tc_wd[51]  = tc_wd[51];
    assign \tc_wd[50]  = tc_wd[50];
    assign \tc_wd[49]  = tc_wd[49];
    assign \tc_wd[48]  = tc_wd[48];
    assign \tc_wd[47]  = tc_wd[47];
    assign \tc_wd[46]  = tc_wd[46];
    assign \tc_wd[45]  = tc_wd[45];
    assign \tc_wd[44]  = tc_wd[44];
    assign \tc_wd[43]  = tc_wd[43];
    assign \tc_wd[40]  = tc_wd[40];
    assign \tc_wd[39]  = tc_wd[39];
    assign \tc_wd[38]  = tc_wd[38];
    assign \tc_wd[36]  = tc_wd[36];
    assign \tc_wd[32]  = tc_wd[32];
    assign \tc_a[60]  = tc_a[60];
    assign \tc_a[58]  = tc_a[58];
    assign ts_i[2] = 1'b0;
    assign ts_i[1] = 1'b0;
    assign ts_i[0] = 1'b0;
    assign adr_i[28] = \tc_a[60] ;
    assign adr_i[26] = \tc_a[58] ;
    assign dat_i[31] = \tc_wd[63] ;
    assign dat_i[30] = \tc_wd[62] ;
    assign dat_i[29] = \tc_wd[61] ;
    assign dat_i[28] = \tc_wd[60] ;
    assign dat_i[27] = \tc_wd[59] ;
    assign dat_i[26] = \tc_wd[58] ;
    assign dat_i[24] = \tc_wd[56] ;
    assign dat_i[23] = \tc_wd[55] ;
    assign dat_i[22] = \tc_wd[54] ;
    assign dat_i[21] = \tc_wd[53] ;
    assign dat_i[20] = \tc_wd[52] ;
    assign dat_i[19] = \tc_wd[51] ;
    assign dat_i[18] = \tc_wd[50] ;
    assign dat_i[17] = \tc_wd[49] ;
    assign dat_i[16] = \tc_wd[48] ;
    assign dat_i[15] = \tc_wd[47] ;
    assign dat_i[14] = \tc_wd[46] ;
    assign dat_i[13] = \tc_wd[45] ;
    assign dat_i[12] = \tc_wd[44] ;
    assign dat_i[11] = \tc_wd[43] ;
    assign dat_i[8] = \tc_wd[40] ;
    assign dat_i[7] = \tc_wd[39] ;
    assign dat_i[6] = \tc_wd[38] ;
    assign dat_i[4] = \tc_wd[36] ;
    assign dat_i[0] = \tc_wd[32] ;
    assign prd_i = 1'b0;
    assign sel_i[3] = \sel_i[2] ;
    assign sel_i[2] = \sel_i[2] ;
    assign sel_i[0] = 1'b1;
    assign tc_ack = ack_in;
    assign ack_out = tr_ack;
    sr2dr_word_8 Urd ( .i(dat_o), .req(n1), .h(tr_rd[63:32]), .l(tr_rd[31:0])
         );
    inv_1 U3 ( .x(n334), .a(tc_a[7]) );
    inv_1 U5 ( .x(n311), .a(tc_a[21]) );
    and2_1 U6 ( .x(n129), .a(n309), .b(n310) );
    inv_1 U7 ( .x(n309), .a(tc_a[6]) );
    inv_1 U9 ( .x(n315), .a(tc_itag[4]) );
    nand2_1 U10 ( .x(n348), .a(n349), .b(n350) );
    inv_1 U11 ( .x(n349), .a(tc_a[12]) );
    inv_1 U12 ( .x(n456), .a(n348) );
    inv_1 U13 ( .x(n336), .a(tc_a[30]) );
    inv_1 U14 ( .x(n457), .a(n345) );
    inv_1 U15 ( .x(n303), .a(tc_a[8]) );
    nand3_1 U16 ( .x(n505), .a(n193), .b(n476), .c(n479) );
    inv_1 U17 ( .x(n229), .a(tc_wd[5]) );
    inv_1 U18 ( .x(n226), .a(tc_wd[3]) );
    inv_1 U19 ( .x(n257), .a(tc_wd[16]) );
    inv_1 U20 ( .x(n263), .a(tc_wd[21]) );
    inv_1 U21 ( .x(n260), .a(tc_wd[19]) );
    nand2_1 U22 ( .x(n268), .a(n269), .b(n270) );
    inv_1 U23 ( .x(n269), .a(tc_wd[23]) );
    inv_1 U24 ( .x(n270), .a(\tc_wd[55] ) );
    nand2_1 U25 ( .x(n265), .a(n266), .b(n267) );
    inv_1 U26 ( .x(n266), .a(tc_wd[20]) );
    inv_1 U27 ( .x(n277), .a(tc_wd[27]) );
    inv_1 U28 ( .x(n252), .a(\tc_wd[47] ) );
    nand2_1 U29 ( .x(n248), .a(n249), .b(n250) );
    inv_1 U30 ( .x(n249), .a(tc_wd[12]) );
    nand2_1 U31 ( .x(n245), .a(n246), .b(n247) );
    inv_1 U32 ( .x(n246), .a(tc_wd[13]) );
    inv_1 U33 ( .x(n247), .a(\tc_wd[45] ) );
    nand2_1 U34 ( .x(n242), .a(n243), .b(n244) );
    inv_1 U35 ( .x(n243), .a(tc_wd[11]) );
    nand2_1 U36 ( .x(n222), .a(n223), .b(n224) );
    inv_1 U37 ( .x(n223), .a(tc_wd[0]) );
    inv_1 U38 ( .x(n220), .a(tc_wd[1]) );
    nand2_1 U39 ( .x(n234), .a(n235), .b(n236) );
    inv_1 U40 ( .x(n235), .a(tc_wd[7]) );
    nand2_1 U41 ( .x(n231), .a(n232), .b(n233) );
    inv_1 U42 ( .x(n232), .a(tc_wd[4]) );
    nand2_1 U43 ( .x(n205), .a(n206), .b(n207) );
    inv_1 U44 ( .x(n206), .a(tc_wd[18]) );
    inv_1 U45 ( .x(n203), .a(tc_wd[10]) );
    nand2_1 U46 ( .x(n199), .a(n200), .b(n201) );
    inv_1 U47 ( .x(n200), .a(tc_wd[6]) );
    inv_1 U48 ( .x(n197), .a(tc_wd[2]) );
    inv_1 U49 ( .x(n218), .a(\tc_wd[46] ) );
    nand2_1 U50 ( .x(n214), .a(n215), .b(n216) );
    inv_1 U51 ( .x(n215), .a(tc_wd[30]) );
    nand2_1 U52 ( .x(n211), .a(n212), .b(n213) );
    inv_1 U53 ( .x(n213), .a(\tc_wd[58] ) );
    nand2_1 U54 ( .x(n208), .a(n209), .b(n210) );
    inv_1 U55 ( .x(n209), .a(tc_wd[22]) );
    inv_1 U56 ( .x(n374), .a(tc_rnw[0]) );
    inv_1 U57 ( .x(n375), .a(tc_rnw[1]) );
    inv_1 U58 ( .x(n368), .a(tc_a[18]) );
    inv_1 U59 ( .x(n244), .a(\tc_wd[43] ) );
    inv_1 U60 ( .x(n251), .a(tc_wd[15]) );
    inv_1 U61 ( .x(n250), .a(\tc_wd[44] ) );
    inv_1 U62 ( .x(n280), .a(tc_wd[29]) );
    inv_1 U63 ( .x(n267), .a(\tc_wd[52] ) );
    inv_1 U64 ( .x(n274), .a(tc_wd[24]) );
    inv_1 U65 ( .x(n271), .a(tc_wd[25]) );
    inv_1 U66 ( .x(n212), .a(tc_wd[26]) );
    inv_1 U67 ( .x(n210), .a(\tc_wd[54] ) );
    inv_1 U68 ( .x(n216), .a(\tc_wd[62] ) );
    inv_1 U69 ( .x(n201), .a(\tc_wd[38] ) );
    inv_1 U70 ( .x(n427), .a(n196) );
    inv_1 U71 ( .x(n207), .a(\tc_wd[50] ) );
    inv_1 U72 ( .x(n424), .a(n202) );
    inv_1 U73 ( .x(n236), .a(\tc_wd[39] ) );
    inv_1 U74 ( .x(n233), .a(\tc_wd[36] ) );
    inv_1 U75 ( .x(n240), .a(tc_wd[8]) );
    inv_1 U76 ( .x(n237), .a(tc_wd[9]) );
    inv_1 U77 ( .x(n224), .a(\tc_wd[32] ) );
    inv_1 U78 ( .x(n413), .a(n219) );
    nand2_1 U79 ( .x(n421), .a(n418), .b(n416) );
    nand2_1 U80 ( .x(n428), .a(n425), .b(n422) );
    nand2_1 U81 ( .x(n414), .a(n411), .b(n408) );
    inv_1 U82 ( .x(n238), .a(tc_wd[41]) );
    inv_1 U83 ( .x(n272), .a(tc_wd[57]) );
    inv_1 U84 ( .x(n350), .a(tc_a[44]) );
    inv_1 U85 ( .x(n351), .a(tc_a[43]) );
    inv_1 U86 ( .x(n366), .a(tc_a[41]) );
    inv_1 U87 ( .x(n335), .a(tc_a[39]) );
    inv_1 U88 ( .x(n310), .a(tc_a[38]) );
    inv_1 U89 ( .x(n355), .a(tc_a[52]) );
    and3_1 U90 ( .x(tc_ok), .a(n531), .b(n532), .c(respond) );
    and2_1 U91 ( .x(tc_slow), .a(respond), .b(acc_o) );
    inv_1 U94 ( .x(n313), .a(tc_itag[5]) );
    and2_1 U95 ( .x(n121), .a(n334), .b(n335) );
    and2_1 U96 ( .x(n122), .a(n359), .b(n360) );
    and2_1 U97 ( .x(n123), .a(n336), .b(n337) );
    and2_1 U98 ( .x(n124), .a(n237), .b(n238) );
    and2_1 U99 ( .x(n125), .a(n251), .b(n252) );
    and2_1 U100 ( .x(n126), .a(n271), .b(n272) );
    and2_1 U101 ( .x(n127), .a(n217), .b(n218) );
    and2_1 U102 ( .x(n128), .a(n311), .b(n312) );
    nor2_1 U103 ( .x(n130), .a(tc_size[3]), .b(tc_size[2]) );
    nand2i_1 U105 ( .x(n284), .a(tc_wd[31]), .b(n285) );
    oa22_1 U106 ( .x(n449), .a(tc_a[27]), .b(tc_a[59]), .c(tc_a[54]), .d(tc_a
        [22]) );
    inv_1 U107 ( .x(n359), .a(tc_a[27]) );
    inv_1 U108 ( .x(n360), .a(tc_a[59]) );
    nand2i_1 U109 ( .x(n282), .a(tc_wd[28]), .b(n283) );
    nor2_1 U110 ( .x(n479), .a(tc_itag[0]), .b(tc_itag[5]) );
    nand4_1 U112 ( .x(n380), .a(n279), .b(n276), .c(n284), .d(n282) );
    aoi21_1 U113 ( .x(n425), .a(n200), .b(n201), .c(n427) );
    oa22_1 U114 ( .x(n397), .a(tc_wd[13]), .b(\tc_wd[45] ), .c(tc_wd[11]), .d(
        \tc_wd[43] ) );
    nor2_1 U115 ( .x(n454), .a(tc_a[20]), .b(tc_a[52]) );
    aoi21_1 U116 ( .x(n422), .a(n206), .b(n207), .c(n424) );
    oa22_1 U117 ( .x(n418), .a(tc_wd[26]), .b(\tc_wd[58] ), .c(tc_wd[22]), .d(
        \tc_wd[54] ) );
    oa22_1 U118 ( .x(n416), .a(tc_wd[14]), .b(\tc_wd[46] ), .c(tc_wd[30]), .d(
        \tc_wd[62] ) );
    inv_1 U119 ( .x(n217), .a(tc_wd[14]) );
    aoi22_1 U120 ( .x(n463), .a(n336), .b(n337), .c(n334), .d(n335) );
    nor2_1 U121 ( .x(n453), .a(tc_a[11]), .b(tc_a[43]) );
    oa22_1 U122 ( .x(n395), .a(tc_wd[15]), .b(\tc_wd[47] ), .c(tc_wd[12]), .d(
        \tc_wd[44] ) );
    oa22_1 U123 ( .x(n404), .a(tc_wd[7]), .b(\tc_wd[39] ), .c(tc_wd[4]), .d(
        \tc_wd[36] ) );
    oa22_1 U124 ( .x(n383), .a(tc_wd[23]), .b(\tc_wd[55] ), .c(tc_wd[20]), .d(
        \tc_wd[52] ) );
    aoi21_1 U125 ( .x(n411), .a(n223), .b(n224), .c(n413) );
    nor2_1 U126 ( .x(n443), .a(tc_a[49]), .b(tc_a[17]) );
    aoi22_1 U127 ( .x(n477), .a(n311), .b(n312), .c(n309), .d(n310) );
    oa21_1 U128 ( .x(n455), .a(tc_a[12]), .b(tc_a[44]), .c(n345) );
    inv_1 U129 ( .x(dat_i[5]), .a(n230) );
    inv_1 U130 ( .x(dat_i[9]), .a(n238) );
    inv_1 U131 ( .x(dat_i[25]), .a(n272) );
    buf_1 U132 ( .x(\sel_i[2] ), .a(tc_size[3]) );
    buf_1 U133 ( .x(adr_i[16]), .a(tc_a[48]) );
    nor2_1 U134 ( .x(n135), .a(tc_a[14]), .b(tc_a[46]) );
    inv_1 U135 ( .x(n305), .a(tc_a[46]) );
    inv_1 U136 ( .x(n487), .a(n302) );
    nand2i_1 U137 ( .x(n445), .a(n446), .b(n442) );
    nor2_1 U138 ( .x(n136), .a(tc_a[29]), .b(tc_a[61]) );
    inv_1 U139 ( .x(n320), .a(tc_a[61]) );
    nand2_1 U140 ( .x(n400), .a(n397), .b(n395) );
    inv_1 U141 ( .x(n137), .a(n340) );
    inv_1 U142 ( .x(dat_i[2]), .a(n198) );
    nand2_1 U143 ( .x(n386), .a(n383), .b(n381) );
    nand3i_1 U144 ( .x(n478), .a(n479), .b(n477), .c(n475) );
    nand2_1 U145 ( .x(n407), .a(n404), .b(n402) );
    inv_1 U146 ( .x(dat_i[10]), .a(n204) );
    inv_1 U147 ( .x(dat_i[1]), .a(n221) );
    nor2_1 U148 ( .x(n141), .a(tc_a[3]), .b(tc_a[35]) );
    inv_1 U149 ( .x(n321), .a(tc_a[35]) );
    nor2_1 U151 ( .x(n483), .a(n484), .b(n485) );
    nor2_1 U152 ( .x(n480), .a(n474), .b(n478) );
    inv_1 U153 ( .x(dat_i[3]), .a(n227) );
    nor2_1 U154 ( .x(n188), .a(n517), .b(n525) );
    nand2_1 U155 ( .x(n180), .a(n401), .b(n387) );
    nor2_1 U156 ( .x(n401), .a(n394), .b(n400) );
    nor2_1 U157 ( .x(n387), .a(n380), .b(n386) );
    nor2_1 U158 ( .x(n481), .a(n482), .b(n135) );
    nor2_1 U159 ( .x(n491), .a(n195), .b(n492) );
    nor2_1 U160 ( .x(n195), .a(tc_size[1]), .b(tc_size[3]) );
    inv_1 U161 ( .x(adr_i[18]), .a(n369) );
    nand2_1 U162 ( .x(n181), .a(n429), .b(n415) );
    nor2_1 U163 ( .x(n429), .a(n421), .b(n428) );
    nor2_1 U164 ( .x(n415), .a(n407), .b(n414) );
    inv_1 U165 ( .x(adr_i[0]), .a(n324) );
    inv_1 U166 ( .x(n324), .a(tc_a[32]) );
    inv_1 U167 ( .x(sel_i[1]), .a(n130) );
    inv_1 U168 ( .x(st_i[2]), .a(n343) );
    inv_1 U169 ( .x(adr_i[9]), .a(n366) );
    inv_1 U170 ( .x(adr_i[24]), .a(n363) );
    inv_1 U171 ( .x(adr_i[19]), .a(n319) );
    inv_1 U172 ( .x(n319), .a(tc_a[51]) );
    inv_1 U173 ( .x(n369), .a(tc_a[50]) );
    inv_1 U174 ( .x(st_i[3]), .a(n344) );
    inv_1 U175 ( .x(adr_i[13]), .a(n354) );
    inv_1 U176 ( .x(adr_i[12]), .a(n350) );
    inv_1 U177 ( .x(adr_i[8]), .a(n304) );
    inv_1 U178 ( .x(n304), .a(tc_a[40]) );
    inv_1 U179 ( .x(adr_i[2]), .a(n330) );
    buf_1 U180 ( .x(adr_i[17]), .a(tc_a[49]) );
    nand2_1 U181 ( .x(n497), .a(n496), .b(n130) );
    inv_1 U182 ( .x(adr_i[10]), .a(n291) );
    and2_1 U183 ( .x(n438), .a(n373), .b(n367) );
    inv_1 U184 ( .x(n439), .a(n373) );
    inv_1 U185 ( .x(n440), .a(n367) );
    inv_1 U186 ( .x(adr_i[20]), .a(n355) );
    inv_1 U187 ( .x(adr_i[27]), .a(n360) );
    inv_1 U188 ( .x(adr_i[4]), .a(n333) );
    inv_1 U189 ( .x(adr_i[25]), .a(n308) );
    inv_1 U190 ( .x(adr_i[30]), .a(n337) );
    inv_1 U191 ( .x(adr_i[31]), .a(n297) );
    inv_1 U192 ( .x(n297), .a(tc_a[63]) );
    inv_1 U193 ( .x(adr_i[15]), .a(n347) );
    inv_1 U194 ( .x(adr_i[11]), .a(n351) );
    inv_1 U195 ( .x(adr_i[1]), .a(n301) );
    inv_1 U196 ( .x(n301), .a(tc_a[33]) );
    nand2_1 U197 ( .x(n503), .a(n499), .b(n502) );
    nor2_1 U198 ( .x(n499), .a(n497), .b(n498) );
    inv_1 U199 ( .x(adr_i[21]), .a(n312) );
    inv_1 U200 ( .x(n312), .a(tc_a[53]) );
    inv_1 U201 ( .x(seq_i), .a(n288) );
    inv_1 U202 ( .x(adr_i[5]), .a(n327) );
    inv_1 U203 ( .x(st_i[4]), .a(n316) );
    inv_1 U204 ( .x(n316), .a(tc_itag[9]) );
    inv_1 U205 ( .x(st_i[1]), .a(n298) );
    inv_1 U206 ( .x(adr_i[23]), .a(n294) );
    inv_1 U207 ( .x(adr_i[22]), .a(n358) );
    nand2_1 U208 ( .x(complb0), .a(n188), .b(n189) );
    nor2_1 U209 ( .x(n189), .a(n503), .b(n510) );
    inv_1 U210 ( .x(adr_i[29]), .a(n320) );
    inv_1 U211 ( .x(adr_i[7]), .a(n335) );
    inv_1 U212 ( .x(adr_i[14]), .a(n305) );
    inv_1 U213 ( .x(adr_i[6]), .a(n310) );
    inv_1 U214 ( .x(st_i[0]), .a(n313) );
    inv_1 U215 ( .x(adr_i[3]), .a(n321) );
    nand3_1 U218 ( .x(n507), .a(n192), .b(n136), .c(n473) );
    nand2_1 U219 ( .x(n508), .a(n471), .b(n141) );
    nor2_1 U220 ( .x(n488), .a(n489), .b(n490) );
    nand4_1 U222 ( .x(complw0), .a(n182), .b(n183), .c(n184), .d(n185) );
    nor2_1 U223 ( .x(n192), .a(\tc_a[58] ), .b(tc_a[26]) );
    nor2_1 U224 ( .x(n193), .a(tc_a[48]), .b(tc_a[16]) );
    nand2_1 U225 ( .x(n364), .a(n365), .b(n366) );
    nand2_1 U226 ( .x(n394), .a(n391), .b(n388) );
    nand4_1 U227 ( .x(n430), .a(n423), .b(n424), .c(n426), .d(n427) );
    nand4_1 U228 ( .x(n431), .a(n127), .b(n417), .c(n419), .d(n420) );
    nor2_1 U229 ( .x(n185), .a(n430), .b(n431) );
    nand4_1 U230 ( .x(n432), .a(n409), .b(n410), .c(n412), .d(n413) );
    nand4_1 U231 ( .x(n433), .a(n403), .b(n124), .c(n405), .d(n406) );
    nor2_1 U232 ( .x(n184), .a(n432), .b(n433) );
    nand4_1 U233 ( .x(n434), .a(n125), .b(n396), .c(n398), .d(n399) );
    nand4_1 U234 ( .x(n435), .a(n389), .b(n390), .c(n392), .d(n393) );
    nor2_1 U235 ( .x(n183), .a(n434), .b(n435) );
    nand4_1 U236 ( .x(n436), .a(n382), .b(n126), .c(n384), .d(n385) );
    nand4_1 U237 ( .x(n437), .a(n376), .b(n377), .c(n378), .d(n379) );
    nor2_1 U238 ( .x(n182), .a(n436), .b(n437) );
    nand2_1 U239 ( .x(n441), .a(n438), .b(n370) );
    nor2_1 U240 ( .x(n442), .a(n443), .b(n444) );
    nor3_1 U241 ( .x(n470), .a(n471), .b(n136), .c(n141) );
    nor3_1 U242 ( .x(n472), .a(n473), .b(n192), .c(n193) );
    nand2_1 U243 ( .x(n474), .a(n472), .b(n470) );
    nor2_1 U244 ( .x(n475), .a(n476), .b(n194) );
    nand3i_1 U245 ( .x(n486), .a(n487), .b(n481), .c(n483) );
    nand3i_1 U246 ( .x(n493), .a(n494), .b(n488), .c(n491) );
    nor2_1 U247 ( .x(n495), .a(n493), .b(n486) );
    nand2_1 U248 ( .x(n191), .a(n495), .b(n480) );
    nand3_1 U249 ( .x(n498), .a(n489), .b(n492), .c(n490) );
    nand3_1 U250 ( .x(n500), .a(n485), .b(n494), .c(n484) );
    nand2_1 U251 ( .x(n501), .a(n135), .b(n487) );
    nor2_1 U252 ( .x(n502), .a(n500), .b(n501) );
    nand3_1 U253 ( .x(n504), .a(n128), .b(n482), .c(n129) );
    nor2_1 U254 ( .x(n506), .a(n504), .b(n505) );
    nor2_1 U255 ( .x(n509), .a(n507), .b(n508) );
    nand2_1 U256 ( .x(n510), .a(n509), .b(n506) );
    nand3_1 U257 ( .x(n511), .a(n465), .b(n466), .c(n468) );
    nand3_1 U258 ( .x(n512), .a(n123), .b(n121), .c(n460) );
    nor2_1 U259 ( .x(n513), .a(n511), .b(n512) );
    nand3_1 U260 ( .x(n514), .a(n462), .b(n459), .c(n457) );
    nand2_1 U261 ( .x(n515), .a(n453), .b(n456) );
    nor2_1 U262 ( .x(n516), .a(n514), .b(n515) );
    nand2_1 U263 ( .x(n517), .a(n516), .b(n513) );
    nand2_1 U264 ( .x(n518), .a(n454), .b(n452) );
    nor2i_1 U265 ( .x(n519), .a(n450), .b(n518) );
    nand2_1 U266 ( .x(n520), .a(n444), .b(n122) );
    nor2i_1 U267 ( .x(n522), .a(n446), .b(n521) );
    nand2_1 U268 ( .x(n523), .a(n439), .b(n524) );
    inv_1 U270 ( .x(n365), .a(tc_a[9]) );
    inv_1 U271 ( .x(n371), .a(\tc_a[60] ) );
    inv_1 U272 ( .x(n446), .a(n364) );
    nor2_1 U273 ( .x(complb1), .a(n190), .b(n191) );
    nor2_1 U274 ( .x(complw1), .a(n180), .b(n181) );
    nand3i_1 U276 ( .x(n190), .a(n441), .b(n447), .c(n469) );
    and4_1 U277 ( .x(n5), .a(n3), .b(n4), .c(n519), .d(n522) );
    inv_1 U216 ( .x(n3), .a(n520) );
    inv_1 U217 ( .x(n4), .a(n523) );
    inv_1 U428 ( .x(n525), .a(n5) );
    nor2_1 U278 ( .x(n447), .a(n448), .b(n445) );
    nor2_1 U279 ( .x(n469), .a(n467), .b(n461) );
    nand2_1 U280 ( .x(n370), .a(n371), .b(n372) );
    nand3i_1 U281 ( .x(n448), .a(n454), .b(n449), .c(n451) );
    nand3i_1 U282 ( .x(n461), .a(n462), .b(n455), .c(n458) );
    nand3i_1 U283 ( .x(n467), .a(n468), .b(n463), .c(n464) );
    inv_1 U284 ( .x(n382), .a(n273) );
    inv_1 U285 ( .x(n384), .a(n268) );
    inv_1 U286 ( .x(n385), .a(n265) );
    inv_1 U287 ( .x(n376), .a(n284) );
    inv_1 U288 ( .x(n377), .a(n282) );
    inv_1 U289 ( .x(n378), .a(n279) );
    inv_1 U290 ( .x(n379), .a(n276) );
    inv_1 U291 ( .x(n396), .a(n248) );
    inv_1 U292 ( .x(n398), .a(n245) );
    inv_1 U293 ( .x(n399), .a(n242) );
    inv_1 U294 ( .x(n389), .a(n262) );
    inv_1 U295 ( .x(n390), .a(n259) );
    inv_1 U296 ( .x(n392), .a(n256) );
    inv_1 U297 ( .x(n393), .a(n253) );
    inv_1 U298 ( .x(n409), .a(n228) );
    inv_1 U299 ( .x(n410), .a(n225) );
    inv_1 U300 ( .x(n412), .a(n222) );
    inv_1 U301 ( .x(n403), .a(n239) );
    inv_1 U302 ( .x(n405), .a(n234) );
    inv_1 U303 ( .x(n406), .a(n231) );
    inv_1 U304 ( .x(n423), .a(n205) );
    inv_1 U305 ( .x(n426), .a(n199) );
    inv_1 U306 ( .x(n417), .a(n214) );
    inv_1 U307 ( .x(n419), .a(n211) );
    inv_1 U308 ( .x(n420), .a(n208) );
    inv_1 U309 ( .x(n444), .a(n361) );
    inv_1 U310 ( .x(n524), .a(n370) );
    inv_1 U311 ( .x(n450), .a(n356) );
    nand2_1 U312 ( .x(n521), .a(n443), .b(n440) );
    inv_1 U313 ( .x(n372), .a(tc_a[28]) );
    nor2_1 U314 ( .x(n451), .a(n452), .b(n453) );
    nor2_1 U315 ( .x(n458), .a(n459), .b(n460) );
    inv_1 U316 ( .x(n468), .a(n331) );
    nor2_1 U317 ( .x(n464), .a(n465), .b(n466) );
    inv_1 U318 ( .x(n494), .a(n295) );
    nand2_1 U319 ( .x(n273), .a(n274), .b(n275) );
    nand2_1 U320 ( .x(n279), .a(n280), .b(n281) );
    nand2_1 U321 ( .x(n276), .a(n277), .b(n278) );
    nand2_1 U322 ( .x(n262), .a(n263), .b(n264) );
    nand2_1 U323 ( .x(n259), .a(n260), .b(n261) );
    nand2_1 U324 ( .x(n256), .a(n257), .b(n258) );
    nand2_1 U325 ( .x(n253), .a(n254), .b(n255) );
    nand2_1 U326 ( .x(n228), .a(n229), .b(n230) );
    nand2_1 U327 ( .x(n225), .a(n226), .b(n227) );
    nand2_1 U328 ( .x(n219), .a(n220), .b(n221) );
    nand2_1 U329 ( .x(n239), .a(n240), .b(n241) );
    nand2_1 U330 ( .x(n202), .a(n203), .b(n204) );
    nand2_1 U331 ( .x(n196), .a(n197), .b(n198) );
    nor2_1 U332 ( .x(n391), .a(n392), .b(n393) );
    nor2_1 U333 ( .x(n388), .a(n389), .b(n390) );
    nor2_1 U334 ( .x(n381), .a(n382), .b(n126) );
    nor2_1 U335 ( .x(n402), .a(n403), .b(n124) );
    nor2_1 U336 ( .x(n408), .a(n409), .b(n410) );
    inv_1 U337 ( .x(n459), .a(n341) );
    inv_1 U338 ( .x(n465), .a(n328) );
    inv_1 U339 ( .x(n466), .a(n325) );
    inv_1 U340 ( .x(n460), .a(n338) );
    nand2_1 U341 ( .x(n361), .a(n362), .b(n363) );
    nand2_1 U342 ( .x(n373), .a(n374), .b(n375) );
    nand2_1 U343 ( .x(n356), .a(n358), .b(n357) );
    inv_1 U344 ( .x(n452), .a(n352) );
    inv_1 U345 ( .x(n484), .a(n299) );
    inv_1 U346 ( .x(n489), .a(n289) );
    inv_1 U347 ( .x(n492), .a(n286) );
    inv_1 U348 ( .x(n490), .a(n292) );
    inv_1 U349 ( .x(n473), .a(n317) );
    inv_1 U350 ( .x(n471), .a(n322) );
    inv_1 U351 ( .x(n482), .a(n306) );
    inv_1 U352 ( .x(n476), .a(n314) );
    nand2_1 U353 ( .x(n367), .a(n368), .b(n369) );
    nand2_1 U354 ( .x(n331), .a(n332), .b(n333) );
    nand2_1 U355 ( .x(n302), .a(n303), .b(n304) );
    nand2_1 U356 ( .x(n295), .a(n296), .b(n297) );
    inv_1 U357 ( .x(n275), .a(\tc_wd[56] ) );
    inv_1 U358 ( .x(n285), .a(\tc_wd[63] ) );
    inv_1 U359 ( .x(n283), .a(\tc_wd[60] ) );
    inv_1 U360 ( .x(n281), .a(\tc_wd[61] ) );
    inv_1 U361 ( .x(n278), .a(\tc_wd[59] ) );
    inv_1 U362 ( .x(n264), .a(\tc_wd[53] ) );
    inv_1 U363 ( .x(n261), .a(\tc_wd[51] ) );
    inv_1 U364 ( .x(n258), .a(\tc_wd[48] ) );
    inv_1 U365 ( .x(n254), .a(tc_wd[17]) );
    inv_1 U366 ( .x(n255), .a(\tc_wd[49] ) );
    inv_1 U367 ( .x(n230), .a(tc_wd[37]) );
    inv_1 U368 ( .x(n227), .a(tc_wd[35]) );
    inv_1 U369 ( .x(n221), .a(tc_wd[33]) );
    inv_1 U370 ( .x(n241), .a(\tc_wd[40] ) );
    inv_1 U371 ( .x(n204), .a(tc_wd[42]) );
    inv_1 U372 ( .x(n198), .a(tc_wd[34]) );
    nand2_1 U373 ( .x(n341), .a(n342), .b(n343) );
    nand2_1 U374 ( .x(n345), .a(n347), .b(n346) );
    nand2_1 U375 ( .x(n328), .a(n329), .b(n330) );
    nand2_1 U376 ( .x(n325), .a(n326), .b(n327) );
    nand2_1 U377 ( .x(n338), .a(n340), .b(n339) );
    inv_1 U378 ( .x(n362), .a(tc_a[24]) );
    inv_1 U379 ( .x(n363), .a(tc_a[56]) );
    inv_1 U380 ( .x(n357), .a(tc_a[22]) );
    inv_1 U381 ( .x(n358), .a(tc_a[54]) );
    nand2_1 U382 ( .x(n352), .a(n353), .b(n354) );
    nand2_1 U383 ( .x(n299), .a(n300), .b(n301) );
    nand2_1 U384 ( .x(n289), .a(n290), .b(n291) );
    nand2_1 U385 ( .x(n286), .a(n287), .b(n288) );
    nand2_1 U386 ( .x(n292), .a(n293), .b(n294) );
    nand2_1 U387 ( .x(n317), .a(n318), .b(n319) );
    nand2_1 U388 ( .x(n322), .a(n323), .b(n324) );
    nand2_1 U389 ( .x(n306), .a(n307), .b(n308) );
    nand2_1 U390 ( .x(n314), .a(n315), .b(n316) );
    inv_1 U391 ( .x(n332), .a(tc_a[4]) );
    inv_1 U392 ( .x(n333), .a(tc_a[36]) );
    inv_1 U393 ( .x(n296), .a(tc_a[31]) );
    inv_1 U394 ( .x(n342), .a(tc_itag[2]) );
    inv_1 U395 ( .x(n343), .a(tc_itag[7]) );
    inv_1 U396 ( .x(n346), .a(tc_a[15]) );
    inv_1 U397 ( .x(n347), .a(tc_a[47]) );
    inv_1 U398 ( .x(n329), .a(tc_a[2]) );
    inv_1 U399 ( .x(n330), .a(tc_a[34]) );
    inv_1 U400 ( .x(n326), .a(tc_a[5]) );
    inv_1 U401 ( .x(n327), .a(tc_a[37]) );
    inv_1 U402 ( .x(n337), .a(tc_a[62]) );
    inv_1 U403 ( .x(n339), .a(tc_lock[0]) );
    inv_1 U404 ( .x(n340), .a(tc_lock[1]) );
    inv_1 U405 ( .x(n353), .a(tc_a[13]) );
    inv_1 U406 ( .x(n354), .a(tc_a[45]) );
    inv_1 U407 ( .x(n300), .a(tc_a[1]) );
    inv_1 U408 ( .x(n290), .a(tc_a[10]) );
    inv_1 U409 ( .x(n291), .a(tc_a[42]) );
    inv_1 U410 ( .x(n287), .a(tc_seq[0]) );
    inv_1 U411 ( .x(n288), .a(tc_seq[1]) );
    inv_1 U412 ( .x(n293), .a(tc_a[23]) );
    inv_1 U413 ( .x(n294), .a(tc_a[55]) );
    inv_1 U414 ( .x(n318), .a(tc_a[19]) );
    inv_1 U415 ( .x(n323), .a(tc_a[0]) );
    inv_1 U416 ( .x(n307), .a(tc_a[25]) );
    inv_1 U417 ( .x(n308), .a(tc_a[57]) );
    buf_1 U418 ( .x(we_i), .a(tc_rnw[0]) );
    matched_delay_cp2slave_resp_dmem U419 ( .x(req_out_delayed), .a(req_out)
         );
    and4_1 U420 ( .x(_25_net_), .a(sel_o[0]), .b(sel_o[1]), .c(n529), .d(n530)
         );
    inv_1 U421 ( .x(_24_net_), .a(we_i) );
    and2_1 U422 ( .x(tc_defer), .a(rty_o), .b(respond) );
    and4_1 U423 ( .x(_26_net_), .a(sel_o[0]), .b(sel_o[1]), .c(sel_o[3]), .d(
        sel_o[2]) );
    inv_1 U424 ( .x(n532), .a(acc_o) );
    inv_1 U425 ( .x(n531), .a(rty_o) );
    inv_1 U426 ( .x(n529), .a(sel_o[2]) );
    inv_1 U427 ( .x(n530), .a(sel_o[3]) );
    buf_1 U150 ( .x(n142), .a(req_in_i) );
    matched_delay_cp2slave_comdmem matchDelCom ( .x(req_in), .a(req_in_i) );
    nand2_1 U275 ( .x(req_in_i), .a(n186), .b(n187) );
    inv_1 U221 ( .x(n186), .a(all_w) );
    inv_1 U269 ( .x(n187), .a(all_r) );
    dffp_1 mult_i_reg ( .q(mult_i), .d(n137), .ck(n142) );
    ao222_1 \cg_respond/__tmp99/U1  ( .x(respond), .a(req_out), .b(tc_ack), 
        .c(req_out), .d(respond), .e(tc_ack), .f(respond) );
    oa21_1 \cg_all_r/__tmp99/U1  ( .x(all_r), .a(tc_rnw[1]), .b(all_r), .c(
        comp_basic) );
    ao31_1 \cg_all_w/__tmp99/aoi  ( .x(\cg_all_w/__tmp99/loop ), .a(comp_basic
        ), .b(comp_wd), .c(we_i), .d(all_w) );
    oa21_1 \cg_all_w/__tmp99/outGate  ( .x(all_w), .a(comp_basic), .b(comp_wd), 
        .c(\cg_all_w/__tmp99/loop ) );
    ao222_1 \cg_wd/__tmp99/U1  ( .x(comp_wd), .a(complw0), .b(complw1), .c(
        complw0), .d(comp_wd), .e(complw1), .f(comp_wd) );
    ao222_1 \cg_basic/__tmp99/U1  ( .x(comp_basic), .a(complb0), .b(complb1), 
        .c(complb0), .d(comp_basic), .e(complb1), .f(comp_basic) );
    inv_1 \Usze1/Uii  ( .x(\Usze1/ni ), .a(_26_net_) );
    inv_1 \Usze1/Uih  ( .x(\Usze1/nh ), .a(tr_size[3]) );
    inv_1 \Usze1/Uil  ( .x(\Usze1/nl ), .a(tr_size[1]) );
    ao23_1 \Usze1/Ucl/U1/U1  ( .x(tr_size[1]), .a(n2), .b(tr_size[1]), .c(n1), 
        .d(\Usze1/ni ), .e(\Usze1/nh ) );
    ao23_1 \Usze1/Uch/U1/U1  ( .x(tr_size[3]), .a(n1), .b(tr_size[3]), .c(n1), 
        .d(_26_net_), .e(\Usze1/nl ) );
    inv_1 \Usze0/Uii  ( .x(\Usze0/ni ), .a(_25_net_) );
    inv_1 \Usze0/Uih  ( .x(\Usze0/nh ), .a(tr_size[2]) );
    inv_1 \Usze0/Uil  ( .x(\Usze0/nl ), .a(tr_size[0]) );
    ao23_1 \Usze0/Ucl/U1/U1  ( .x(tr_size[0]), .a(n2), .b(tr_size[0]), .c(n1), 
        .d(\Usze0/ni ), .e(\Usze0/nh ) );
    ao23_1 \Usze0/Uch/U1/U1  ( .x(tr_size[2]), .a(n2), .b(tr_size[2]), .c(n1), 
        .d(_25_net_), .e(\Usze0/nl ) );
    inv_1 \Urnw/Uii  ( .x(\Urnw/ni ), .a(_24_net_) );
    inv_1 \Urnw/Uih  ( .x(\Urnw/nh ), .a(tr_rnw[1]) );
    inv_1 \Urnw/Uil  ( .x(\Urnw/nl ), .a(tr_rnw[0]) );
    ao23_1 \Urnw/Ucl/U1/U1  ( .x(tr_rnw[0]), .a(n1), .b(tr_rnw[0]), .c(n1), 
        .d(\Urnw/ni ), .e(\Urnw/nh ) );
    ao23_1 \Urnw/Uch/U1/U1  ( .x(tr_rnw[1]), .a(n1), .b(tr_rnw[1]), .c(n1), 
        .d(_24_net_), .e(\Urnw/nl ) );
    inv_1 \Uerr/Uii  ( .x(\Uerr/ni ), .a(err_o) );
    inv_1 \Uerr/Uih  ( .x(\Uerr/nh ), .a(tr_err[1]) );
    inv_1 \Uerr/Uil  ( .x(\Uerr/nl ), .a(tr_err[0]) );
    ao23_1 \Uerr/Ucl/U1/U1  ( .x(tr_err[0]), .a(n1), .b(tr_err[0]), .c(n1), 
        .d(\Uerr/ni ), .e(\Uerr/nh ) );
    ao23_1 \Uerr/Uch/U1/U1  ( .x(tr_err[1]), .a(n1), .b(tr_err[1]), .c(n1), 
        .d(err_o), .e(\Uerr/nl ) );
    inv_0 U1 ( .x(n298), .a(tc_itag[6]) );
    nor2_0 U2 ( .x(n485), .a(tc_itag[1]), .b(tc_itag[6]) );
    inv_0 U4 ( .x(n344), .a(tc_itag[8]) );
    nor2_0 U8 ( .x(n462), .a(tc_itag[3]), .b(tc_itag[8]) );
    nor2_0 U92 ( .x(n496), .a(tc_size[0]), .b(tc_size[1]) );
    nor2_0 U93 ( .x(n194), .a(tc_size[0]), .b(tc_size[2]) );
    buf_16 U104 ( .x(n1), .a(req_out_delayed) );
    buf_16 U111 ( .x(n2), .a(req_out_delayed) );
endmodule


module slave_if_dmem ( nReset, sc_req, sc_we, sc_mult, sc_seq, sc_prd, sc_ts, 
    sc_st, sc_sel, sc_adr, sc_dat, sc_ack, sr_req, sr_err, sr_rty, sr_acc, 
    sr_mult, sr_ts, sr_rt, sr_sel, sr_dat, sr_ack, chaincommand, 
    nchaincommandack, chainresponse, nchainresponseack, e_dp, e_ip, e_tic, 
    r_dp, r_ip, r_tic );
output [2:0] sc_ts;
output [4:0] sc_st;
output [3:0] sc_sel;
output [31:0] sc_adr;
output [31:0] sc_dat;
input  [2:0] sr_ts;
input  [4:0] sr_rt;
input  [3:0] sr_sel;
input  [31:0] sr_dat;
input  [4:0] chaincommand;
output [4:0] chainresponse;
input  [2:0] e_dp;
input  [2:0] e_ip;
input  [2:0] e_tic;
input  [2:0] r_dp;
input  [2:0] r_ip;
input  [2:0] r_tic;
input  nReset, sc_ack, sr_req, sr_err, sr_rty, sr_acc, sr_mult, 
    nchainresponseack;
output sc_req, sc_we, sc_mult, sc_seq, sc_prd, sr_ack, nchaincommandack;
    wire \ct_a[63] , \ct_a[62] , \ct_a[61] , \ct_a[60] , \ct_a[59] , 
        \ct_a[58] , \ct_a[57] , \ct_a[56] , \ct_a[55] , \ct_a[54] , \ct_a[53] , 
        \ct_a[52] , \ct_a[51] , \ct_a[50] , \ct_a[49] , \ct_a[48] , \ct_a[47] , 
        \ct_a[46] , \ct_a[45] , \ct_a[44] , \ct_a[43] , \ct_a[42] , \ct_a[41] , 
        \ct_a[40] , \ct_a[39] , \ct_a[38] , \ct_a[37] , \ct_a[36] , \ct_a[35] , 
        \ct_a[34] , \ct_a[33] , \ct_a[32] , \ct_a[31] , \ct_a[30] , \ct_a[29] , 
        \ct_a[28] , \ct_a[27] , \ct_a[26] , \ct_a[25] , \ct_a[24] , \ct_a[23] , 
        \ct_a[22] , \ct_a[21] , \ct_a[20] , \ct_a[19] , \ct_a[18] , \ct_a[17] , 
        \ct_a[16] , \ct_a[15] , \ct_a[14] , \ct_a[13] , \ct_a[12] , \ct_a[11] , 
        \ct_a[10] , \ct_a[9] , \ct_a[8] , \ct_a[7] , \ct_a[6] , \ct_a[5] , 
        \ct_a[4] , \ct_a[3] , \ct_a[2] , \ct_a[1] , \ct_a[0] , \ct_wd[63] , 
        \ct_wd[62] , \ct_wd[61] , \ct_wd[60] , \ct_wd[59] , \ct_wd[58] , 
        \ct_wd[57] , \ct_wd[56] , \ct_wd[55] , \ct_wd[54] , \ct_wd[53] , 
        \ct_wd[52] , \ct_wd[51] , \ct_wd[50] , \ct_wd[49] , \ct_wd[48] , 
        \ct_wd[47] , \ct_wd[46] , \ct_wd[45] , \ct_wd[44] , \ct_wd[43] , 
        \ct_wd[42] , \ct_wd[41] , \ct_wd[40] , \ct_wd[39] , \ct_wd[38] , 
        \ct_wd[37] , \ct_wd[36] , \ct_wd[35] , \ct_wd[34] , \ct_wd[33] , 
        \ct_wd[32] , \ct_wd[31] , \ct_wd[30] , \ct_wd[29] , \ct_wd[28] , 
        \ct_wd[27] , \ct_wd[26] , \ct_wd[25] , \ct_wd[24] , \ct_wd[23] , 
        \ct_wd[22] , \ct_wd[21] , \ct_wd[20] , \ct_wd[19] , \ct_wd[18] , 
        \ct_wd[17] , \ct_wd[16] , \ct_wd[15] , \ct_wd[14] , \ct_wd[13] , 
        \ct_wd[12] , \ct_wd[11] , \ct_wd[10] , \ct_wd[9] , \ct_wd[8] , 
        \ct_wd[7] , \ct_wd[6] , \ct_wd[5] , \ct_wd[4] , \ct_wd[3] , \ct_wd[2] , 
        \ct_wd[1] , \ct_wd[0] , \ct_rnw[1] , \ct_rnw[0] , \ct_lock[1] , 
        \ct_lock[0] , \ct_seq[1] , \ct_seq[0] , \ct_size[3] , \ct_size[2] , 
        \ct_size[1] , \ct_size[0] , \ct_itag[9] , \ct_itag[8] , \ct_itag[7] , 
        \ct_itag[6] , \ct_itag[5] , \ct_itag[4] , \ct_itag[3] , \ct_itag[2] , 
        \ct_itag[1] , \ct_itag[0] , ct_ack, ct_ok, ct_defer, ct_slow, 
        \rt_rd[63] , \rt_rd[62] , \rt_rd[61] , \rt_rd[60] , \rt_rd[59] , 
        \rt_rd[58] , \rt_rd[57] , \rt_rd[56] , \rt_rd[55] , \rt_rd[54] , 
        \rt_rd[53] , \rt_rd[52] , \rt_rd[51] , \rt_rd[50] , \rt_rd[49] , 
        \rt_rd[48] , \rt_rd[47] , \rt_rd[46] , \rt_rd[45] , \rt_rd[44] , 
        \rt_rd[43] , \rt_rd[42] , \rt_rd[41] , \rt_rd[40] , \rt_rd[39] , 
        \rt_rd[38] , \rt_rd[37] , \rt_rd[36] , \rt_rd[35] , \rt_rd[34] , 
        \rt_rd[33] , \rt_rd[32] , \rt_rd[31] , \rt_rd[30] , \rt_rd[29] , 
        \rt_rd[28] , \rt_rd[27] , \rt_rd[26] , \rt_rd[25] , \rt_rd[24] , 
        \rt_rd[23] , \rt_rd[22] , \rt_rd[21] , \rt_rd[20] , \rt_rd[19] , 
        \rt_rd[18] , \rt_rd[17] , \rt_rd[16] , \rt_rd[15] , \rt_rd[14] , 
        \rt_rd[13] , \rt_rd[12] , \rt_rd[11] , \rt_rd[10] , \rt_rd[9] , 
        \rt_rd[8] , \rt_rd[7] , \rt_rd[6] , \rt_rd[5] , \rt_rd[4] , \rt_rd[3] , 
        \rt_rd[2] , \rt_rd[1] , \rt_rd[0] , \rt_err[1] , \rt_err[0] , rt_ack, 
        \tag_h[4] , \tag_h[3] , \tag_h[2] , \tag_h[1] , \tag_h[0] , \tag_l[4] , 
        \tag_l[3] , \tag_l[2] , \tag_l[1] , \tag_l[0] , \route[4] , \route[1] , 
        \route[0] , nroute_ack, routetx_req, routetx_ack, \eh[1] , \eh[0] , 
        \el[2] , \el[1] , \el[0] , \rh[2] , \rh[1] , \rl[2] , \rl[1] , \rl[0] , 
        reset;
    wire SYNOPSYS_UNCONNECTED_1 , SYNOPSYS_UNCONNECTED_2 , 
	SYNOPSYS_UNCONNECTED_3 , SYNOPSYS_UNCONNECTED_4 , SYNOPSYS_UNCONNECTED_5 ;
    assign sc_prd = 1'b0;
    assign sc_ts[2] = 1'b0;
    assign sc_ts[1] = 1'b0;
    assign sc_ts[0] = 1'b0;
    assign sc_sel[0] = 1'b1;
    target_dmem tg ( .addr({\ct_a[63] , \ct_a[62] , \ct_a[61] , \ct_a[60] , 
        \ct_a[59] , \ct_a[58] , \ct_a[57] , \ct_a[56] , \ct_a[55] , \ct_a[54] , 
        \ct_a[53] , \ct_a[52] , \ct_a[51] , \ct_a[50] , \ct_a[49] , \ct_a[48] , 
        \ct_a[47] , \ct_a[46] , \ct_a[45] , \ct_a[44] , \ct_a[43] , \ct_a[42] , 
        \ct_a[41] , \ct_a[40] , \ct_a[39] , \ct_a[38] , \ct_a[37] , \ct_a[36] , 
        \ct_a[35] , \ct_a[34] , \ct_a[33] , \ct_a[32] , \ct_a[31] , \ct_a[30] , 
        \ct_a[29] , \ct_a[28] , \ct_a[27] , \ct_a[26] , \ct_a[25] , \ct_a[24] , 
        \ct_a[23] , \ct_a[22] , \ct_a[21] , \ct_a[20] , \ct_a[19] , \ct_a[18] , 
        \ct_a[17] , \ct_a[16] , \ct_a[15] , \ct_a[14] , \ct_a[13] , \ct_a[12] , 
        \ct_a[11] , \ct_a[10] , \ct_a[9] , \ct_a[8] , \ct_a[7] , \ct_a[6] , 
        \ct_a[5] , \ct_a[4] , \ct_a[3] , \ct_a[2] , \ct_a[1] , \ct_a[0] }), 
        .chainresponse(chainresponse), .crnw({\ct_rnw[1] , \ct_rnw[0] }), 
        .csize({\ct_size[3] , \ct_size[2] , \ct_size[1] , \ct_size[0] }), 
        .ctag({\ct_itag[9] , \ct_itag[8] , \ct_itag[7] , \ct_itag[6] , 
        \ct_itag[5] , \ct_itag[4] , \ct_itag[3] , \ct_itag[2] , \ct_itag[1] , 
        \ct_itag[0] }), .lock({\ct_lock[1] , \ct_lock[0] }), 
        .nchaincommandack(nchaincommandack), .nrouteack(nroute_ack), .rack(
        rt_ack), .routetxreq(routetx_req), .seq({\ct_seq[1] , \ct_seq[0] }), 
        .tag_h({\tag_h[4] , \tag_h[3] , \tag_h[2] , \tag_h[1] , \tag_h[0] }), 
        .tag_l({\tag_l[4] , \tag_l[3] , \tag_l[2] , \tag_l[1] , \tag_l[0] }), 
        .wd({\ct_wd[63] , \ct_wd[62] , \ct_wd[61] , \ct_wd[60] , \ct_wd[59] , 
        \ct_wd[58] , \ct_wd[57] , \ct_wd[56] , \ct_wd[55] , \ct_wd[54] , 
        \ct_wd[53] , \ct_wd[52] , \ct_wd[51] , \ct_wd[50] , \ct_wd[49] , 
        \ct_wd[48] , \ct_wd[47] , \ct_wd[46] , \ct_wd[45] , \ct_wd[44] , 
        \ct_wd[43] , \ct_wd[42] , \ct_wd[41] , \ct_wd[40] , \ct_wd[39] , 
        \ct_wd[38] , \ct_wd[37] , \ct_wd[36] , \ct_wd[35] , \ct_wd[34] , 
        \ct_wd[33] , \ct_wd[32] , \ct_wd[31] , \ct_wd[30] , \ct_wd[29] , 
        \ct_wd[28] , \ct_wd[27] , \ct_wd[26] , \ct_wd[25] , \ct_wd[24] , 
        \ct_wd[23] , \ct_wd[22] , \ct_wd[21] , \ct_wd[20] , \ct_wd[19] , 
        \ct_wd[18] , \ct_wd[17] , \ct_wd[16] , \ct_wd[15] , \ct_wd[14] , 
        \ct_wd[13] , \ct_wd[12] , \ct_wd[11] , \ct_wd[10] , \ct_wd[9] , 
        \ct_wd[8] , \ct_wd[7] , \ct_wd[6] , \ct_wd[5] , \ct_wd[4] , \ct_wd[3] , 
        \ct_wd[2] , \ct_wd[1] , \ct_wd[0] }), .cack(ct_ack), .cdefer(ct_defer), 
        .chaincommand(chaincommand), .cndefer(ct_slow), .cok(ct_ok), .err({
        \rt_err[1] , \rt_err[0] }), .nReset(nReset), .nchainresponseack(
        nchainresponseack), .rd({\rt_rd[63] , \rt_rd[62] , \rt_rd[61] , 
        \rt_rd[60] , \rt_rd[59] , \rt_rd[58] , \rt_rd[57] , \rt_rd[56] , 
        \rt_rd[55] , \rt_rd[54] , \rt_rd[53] , \rt_rd[52] , \rt_rd[51] , 
        \rt_rd[50] , \rt_rd[49] , \rt_rd[48] , \rt_rd[47] , \rt_rd[46] , 
        \rt_rd[45] , \rt_rd[44] , \rt_rd[43] , \rt_rd[42] , \rt_rd[41] , 
        \rt_rd[40] , \rt_rd[39] , \rt_rd[38] , \rt_rd[37] , \rt_rd[36] , 
        \rt_rd[35] , \rt_rd[34] , \rt_rd[33] , \rt_rd[32] , \rt_rd[31] , 
        \rt_rd[30] , \rt_rd[29] , \rt_rd[28] , \rt_rd[27] , \rt_rd[26] , 
        \rt_rd[25] , \rt_rd[24] , \rt_rd[23] , \rt_rd[22] , \rt_rd[21] , 
        \rt_rd[20] , \rt_rd[19] , \rt_rd[18] , \rt_rd[17] , \rt_rd[16] , 
        \rt_rd[15] , \rt_rd[14] , \rt_rd[13] , \rt_rd[12] , \rt_rd[11] , 
        \rt_rd[10] , \rt_rd[9] , \rt_rd[8] , \rt_rd[7] , \rt_rd[6] , 
        \rt_rd[5] , \rt_rd[4] , \rt_rd[3] , \rt_rd[2] , \rt_rd[1] , \rt_rd[0] 
        }), .route({\route[4] , 1'b0, 1'b0, \route[1] , \route[0] }), 
        .routetxack(routetx_ack) );
    t_adec_dmem dec ( .e_h({SYNOPSYS_UNCONNECTED_1, \eh[1] , \eh[0] }), .e_l({
        \el[2] , \el[1] , \el[0] }), .r_h({\rh[2] , \rh[1] , 
        SYNOPSYS_UNCONNECTED_2}), .r_l({\rl[2] , \rl[1] , \rl[0] }), .e_dp(
        e_dp), .e_ip(e_ip), .e_tic(e_tic), .r_dp(r_dp), .r_ip(r_ip), .r_tic(
        r_tic), .tag_h({\tag_h[4] , \tag_h[3] , \tag_h[2] , \tag_h[1] , 
        \tag_h[0] }), .tag_l({\tag_l[4] , \tag_l[3] , \tag_l[2] , \tag_l[1] , 
        \tag_l[0] }) );
    resp_route_tx_dmem rt ( .o({\route[4] , SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, \route[1] , \route[0] }), .rtxack(routetx_ack), 
        .e_h({1'b0, \eh[1] , \eh[0] }), .e_l({\el[2] , \el[1] , \el[0] }), 
        .noa(nroute_ack), .r_h({\rh[2] , \rh[1] , 1'b0}), .r_l({\rl[2] , 
        \rl[1] , \rl[0] }), .rtxreq(routetx_req) );
    inv_2 U1 ( .x(reset), .a(nReset) );
    cp2slave_dmem chainif2slave ( .tc_seq({\ct_seq[1] , \ct_seq[0] }), 
        .tc_size({\ct_size[3] , \ct_size[2] , \ct_size[1] , \ct_size[0] }), 
        .tc_itag({\ct_itag[9] , \ct_itag[8] , \ct_itag[7] , \ct_itag[6] , 
        \ct_itag[5] , \ct_itag[4] , \ct_itag[3] , \ct_itag[2] , \ct_itag[1] , 
        \ct_itag[0] }), .tc_wd({\ct_wd[63] , \ct_wd[62] , \ct_wd[61] , 
        \ct_wd[60] , \ct_wd[59] , \ct_wd[58] , \ct_wd[57] , \ct_wd[56] , 
        \ct_wd[55] , \ct_wd[54] , \ct_wd[53] , \ct_wd[52] , \ct_wd[51] , 
        \ct_wd[50] , \ct_wd[49] , \ct_wd[48] , \ct_wd[47] , \ct_wd[46] , 
        \ct_wd[45] , \ct_wd[44] , \ct_wd[43] , \ct_wd[42] , \ct_wd[41] , 
        \ct_wd[40] , \ct_wd[39] , \ct_wd[38] , \ct_wd[37] , \ct_wd[36] , 
        \ct_wd[35] , \ct_wd[34] , \ct_wd[33] , \ct_wd[32] , \ct_wd[31] , 
        \ct_wd[30] , \ct_wd[29] , \ct_wd[28] , \ct_wd[27] , \ct_wd[26] , 
        \ct_wd[25] , \ct_wd[24] , \ct_wd[23] , \ct_wd[22] , \ct_wd[21] , 
        \ct_wd[20] , \ct_wd[19] , \ct_wd[18] , \ct_wd[17] , \ct_wd[16] , 
        \ct_wd[15] , \ct_wd[14] , \ct_wd[13] , \ct_wd[12] , \ct_wd[11] , 
        \ct_wd[10] , \ct_wd[9] , \ct_wd[8] , \ct_wd[7] , \ct_wd[6] , 
        \ct_wd[5] , \ct_wd[4] , \ct_wd[3] , \ct_wd[2] , \ct_wd[1] , \ct_wd[0] 
        }), .tc_lock({\ct_lock[1] , \ct_lock[0] }), .tc_a({\ct_a[63] , 
        \ct_a[62] , \ct_a[61] , \ct_a[60] , \ct_a[59] , \ct_a[58] , \ct_a[57] , 
        \ct_a[56] , \ct_a[55] , \ct_a[54] , \ct_a[53] , \ct_a[52] , \ct_a[51] , 
        \ct_a[50] , \ct_a[49] , \ct_a[48] , \ct_a[47] , \ct_a[46] , \ct_a[45] , 
        \ct_a[44] , \ct_a[43] , \ct_a[42] , \ct_a[41] , \ct_a[40] , \ct_a[39] , 
        \ct_a[38] , \ct_a[37] , \ct_a[36] , \ct_a[35] , \ct_a[34] , \ct_a[33] , 
        \ct_a[32] , \ct_a[31] , \ct_a[30] , \ct_a[29] , \ct_a[28] , \ct_a[27] , 
        \ct_a[26] , \ct_a[25] , \ct_a[24] , \ct_a[23] , \ct_a[22] , \ct_a[21] , 
        \ct_a[20] , \ct_a[19] , \ct_a[18] , \ct_a[17] , \ct_a[16] , \ct_a[15] , 
        \ct_a[14] , \ct_a[13] , \ct_a[12] , \ct_a[11] , \ct_a[10] , \ct_a[9] , 
        \ct_a[8] , \ct_a[7] , \ct_a[6] , \ct_a[5] , \ct_a[4] , \ct_a[3] , 
        \ct_a[2] , \ct_a[1] , \ct_a[0] }), .tc_rnw({\ct_rnw[1] , \ct_rnw[0] }), 
        .tc_ok(ct_ok), .tc_defer(ct_defer), .tc_slow(ct_slow), .tc_ack(ct_ack), 
        .req_in(sc_req), .st_i(sc_st), .we_i(sc_we), .mult_i(sc_mult), .adr_i(
        sc_adr), .dat_i(sc_dat), .seq_i(sc_seq), .sel_i({sc_sel[3], sc_sel[2], 
        sc_sel[1], SYNOPSYS_UNCONNECTED_5}), .ack_in(sc_ack), .tr_rd({
        \rt_rd[63] , \rt_rd[62] , \rt_rd[61] , \rt_rd[60] , \rt_rd[59] , 
        \rt_rd[58] , \rt_rd[57] , \rt_rd[56] , \rt_rd[55] , \rt_rd[54] , 
        \rt_rd[53] , \rt_rd[52] , \rt_rd[51] , \rt_rd[50] , \rt_rd[49] , 
        \rt_rd[48] , \rt_rd[47] , \rt_rd[46] , \rt_rd[45] , \rt_rd[44] , 
        \rt_rd[43] , \rt_rd[42] , \rt_rd[41] , \rt_rd[40] , \rt_rd[39] , 
        \rt_rd[38] , \rt_rd[37] , \rt_rd[36] , \rt_rd[35] , \rt_rd[34] , 
        \rt_rd[33] , \rt_rd[32] , \rt_rd[31] , \rt_rd[30] , \rt_rd[29] , 
        \rt_rd[28] , \rt_rd[27] , \rt_rd[26] , \rt_rd[25] , \rt_rd[24] , 
        \rt_rd[23] , \rt_rd[22] , \rt_rd[21] , \rt_rd[20] , \rt_rd[19] , 
        \rt_rd[18] , \rt_rd[17] , \rt_rd[16] , \rt_rd[15] , \rt_rd[14] , 
        \rt_rd[13] , \rt_rd[12] , \rt_rd[11] , \rt_rd[10] , \rt_rd[9] , 
        \rt_rd[8] , \rt_rd[7] , \rt_rd[6] , \rt_rd[5] , \rt_rd[4] , \rt_rd[3] , 
        \rt_rd[2] , \rt_rd[1] , \rt_rd[0] }), .tr_err({\rt_err[1] , 
        \rt_err[0] }), .tr_ack(rt_ack), .req_out(sr_req), .dat_o(sr_dat), 
        .err_o(sr_err), .rty_o(sr_rty), .acc_o(sr_acc), .sel_o(sr_sel), 
        .mult_o(sr_mult), .rt_o(sr_rt), .ack_out(sr_ack), .reset(reset) );
endmodule


module aspida_net_core ( nrst, clk, ip_c_req, ip_c_we, ip_c_mult, ip_c_prd, 
    ip_c_seq, ip_c_ts, ip_c_sel, ip_c_adr, ip_c_dat, ip_c_ack, ip_r_req, 
    ip_r_we, ip_r_err, ip_r_rty, ip_r_acc, ip_r_ts, ip_r_sel, ip_r_dat, 
    ip_r_ack, dp_c_req, dp_c_we, dp_c_mult, dp_c_prd, dp_c_seq, dp_c_ts, 
    dp_c_sel, dp_c_adr, dp_c_dat, dp_c_ack, dp_r_req, dp_r_we, dp_r_err, 
    dp_r_rty, dp_r_acc, dp_r_ts, dp_r_sel, dp_r_dat, dp_r_ack, ei_c_req, 
    ei_c_ack, ei_c_we, ei_c_addr, ei_r_req, ei_r_ack, ei_data_in, ei_data_out, 
    c_BC, c_BC_ack, r_BC, r_BC_ack, wish_we_o, wish_stb_cyc_o, wish_ack_i, 
    wish_adr_o, wish_dat_i, wish_dat_o, dm_c_req, dm_c_we, dm_c_mult, dm_c_seq, 
    dm_c_prd, dm_c_ts, dm_c_st, dm_c_sel, dm_c_adr, dm_c_dat, dm_c_ack, 
    dm_r_req, dm_r_err, dm_r_rty, dm_r_acc, dm_r_mult, dm_r_ts, dm_r_rt, 
    dm_r_sel, dm_r_dat, dm_r_ack, im_c_req, im_c_we, im_c_mult, im_c_seq, 
    im_c_prd, im_c_ts, im_c_st, im_c_sel, im_c_adr, im_c_dat, im_c_ack, 
    im_r_req, im_r_err, im_r_rty, im_r_acc, im_r_mult, im_r_ts, im_r_rt, 
    im_r_sel, im_r_dat, im_r_ack, test_si, test_so, test_se, phi1, phi2, phi3, 
    force_bare );
input  [2:0] ip_c_ts;
input  [3:0] ip_c_sel;
input  [31:0] ip_c_adr;
input  [31:0] ip_c_dat;
output [2:0] ip_r_ts;
output [3:0] ip_r_sel;
output [31:0] ip_r_dat;
input  [2:0] dp_c_ts;
input  [3:0] dp_c_sel;
input  [31:0] dp_c_adr;
input  [31:0] dp_c_dat;
output [2:0] dp_r_ts;
output [3:0] dp_r_sel;
output [31:0] dp_r_dat;
input  [10:0] ei_c_addr;
input  [7:0] ei_data_in;
output [7:0] ei_data_out;
output [4:0] c_BC;
input  [4:0] r_BC;
output [11:0] wish_adr_o;
input  [31:0] wish_dat_i;
output [31:0] wish_dat_o;
output [2:0] dm_c_ts;
output [4:0] dm_c_st;
output [3:0] dm_c_sel;
output [31:0] dm_c_adr;
output [31:0] dm_c_dat;
input  [2:0] dm_r_ts;
input  [4:0] dm_r_rt;
input  [3:0] dm_r_sel;
input  [31:0] dm_r_dat;
output [2:0] im_c_ts;
output [4:0] im_c_st;
output [3:0] im_c_sel;
output [31:0] im_c_adr;
output [31:0] im_c_dat;
input  [2:0] im_r_ts;
input  [4:0] im_r_rt;
input  [3:0] im_r_sel;
input  [31:0] im_r_dat;
input  nrst, clk, ip_c_req, ip_c_we, ip_c_mult, ip_c_prd, ip_c_seq, ip_r_ack, 
    dp_c_req, dp_c_we, dp_c_mult, dp_c_prd, dp_c_seq, dp_r_ack, ei_c_req, 
    ei_c_we, ei_r_ack, c_BC_ack, wish_ack_i, dm_c_ack, dm_r_req, dm_r_err, 
    dm_r_rty, dm_r_acc, dm_r_mult, im_c_ack, im_r_req, im_r_err, im_r_rty, 
    im_r_acc, im_r_mult, test_si, test_se, phi1, phi2, phi3, force_bare;
output ip_c_ack, ip_r_req, ip_r_we, ip_r_err, ip_r_rty, ip_r_acc, dp_c_ack, 
    dp_r_req, dp_r_we, dp_r_err, dp_r_rty, dp_r_acc, ei_c_ack, ei_r_req, 
    r_BC_ack, wish_we_o, wish_stb_cyc_o, dm_c_req, dm_c_we, dm_c_mult, 
    dm_c_seq, dm_c_prd, dm_r_ack, im_c_req, im_c_we, im_c_mult, im_c_seq, 
    im_c_prd, im_r_ack, test_so;
    wire rst, real_c_Iport_ack, c_Iport_ack, \c_Iport[4] , \c_Iport[3] , 
        \c_Iport[2] , \c_Iport[1] , \c_Iport[0] , \r_Iport[4] , \r_Iport[3] , 
        \r_Iport[2] , \r_Iport[1] , \r_Iport[0] , r_Iport_ack, 
        real_c_Dport_ack, c_Dport_ack, \c_Dport[4] , \c_Dport[3] , 
        \c_Dport[2] , \c_Dport[1] , \c_Dport[0] , \r_Dport[4] , \r_Dport[3] , 
        \r_Dport[2] , \r_Dport[1] , \r_Dport[0] , r_Dport_ack, real_c_TIC_ack, 
        c_TIC_ack, tic_c_req, tic_c_we, \tic_c_adr[31] , \tic_c_adr[30] , 
        \tic_c_adr[11] , \tic_c_adr[10] , \tic_c_adr[9] , \tic_c_adr[8] , 
        \tic_c_adr[7] , \tic_c_adr[6] , \tic_c_adr[5] , \tic_c_adr[4] , 
        \tic_c_adr[3] , \tic_c_adr[2] , \tic_c_dat[31] , \tic_c_dat[30] , 
        \tic_c_dat[29] , \tic_c_dat[28] , \tic_c_dat[27] , \tic_c_dat[26] , 
        \tic_c_dat[25] , \tic_c_dat[24] , \tic_c_dat[23] , \tic_c_dat[22] , 
        \tic_c_dat[21] , \tic_c_dat[20] , \tic_c_dat[19] , \tic_c_dat[18] , 
        \tic_c_dat[17] , \tic_c_dat[16] , \tic_c_dat[15] , \tic_c_dat[14] , 
        \tic_c_dat[13] , \tic_c_dat[12] , \tic_c_dat[11] , \tic_c_dat[10] , 
        \tic_c_dat[9] , \tic_c_dat[8] , \tic_c_dat[7] , \tic_c_dat[6] , 
        \tic_c_dat[5] , \tic_c_dat[4] , \tic_c_dat[3] , \tic_c_dat[2] , 
        \tic_c_dat[1] , \tic_c_dat[0] , tic_c_ack, tic_r_req, \tic_r_dat[31] , 
        \tic_r_dat[30] , \tic_r_dat[29] , \tic_r_dat[28] , \tic_r_dat[27] , 
        \tic_r_dat[26] , \tic_r_dat[25] , \tic_r_dat[24] , \tic_r_dat[23] , 
        \tic_r_dat[22] , \tic_r_dat[21] , \tic_r_dat[20] , \tic_r_dat[19] , 
        \tic_r_dat[18] , \tic_r_dat[17] , \tic_r_dat[16] , \tic_r_dat[15] , 
        \tic_r_dat[14] , \tic_r_dat[13] , \tic_r_dat[12] , \tic_r_dat[11] , 
        \tic_r_dat[10] , \tic_r_dat[9] , \tic_r_dat[8] , \tic_r_dat[7] , 
        \tic_r_dat[6] , \tic_r_dat[5] , \tic_r_dat[4] , \tic_r_dat[3] , 
        \tic_r_dat[2] , \tic_r_dat[1] , \tic_r_dat[0] , tic_r_ack, \c_TIC[4] , 
        \c_TIC[3] , \c_TIC[2] , \c_TIC[1] , \c_TIC[0] , \r_TIC[4] , \r_TIC[3] , 
        \r_TIC[2] , \r_TIC[1] , \r_TIC[0] , r_TIC_ack, c_BC_ack_n, c_WB_ack_n, 
        c_WB_ack, c_IMEM_ack_n, c_IMEM_ack, c_DMEM_ack_n, c_DMEM_ack, 
        \c_WB[4] , \c_WB[3] , \c_WB[2] , \c_WB[1] , \c_WB[0] , \c_IMEM[4] , 
        \c_IMEM[3] , \c_IMEM[2] , \c_IMEM[1] , \c_IMEM[0] , \c_DMEM[4] , 
        \c_DMEM[3] , \c_DMEM[2] , \c_DMEM[1] , \c_DMEM[0] , scan_o_cmd, 
        r_Iport_ack_n, r_TIC_ack_n, r_Dport_ack_n, \r_IMEM[4] , \r_IMEM[3] , 
        \r_IMEM[2] , \r_IMEM[1] , \r_IMEM[0] , r_IMEM_ack, \r_DMEM[4] , 
        \r_DMEM[3] , \r_DMEM[2] , \r_DMEM[1] , \r_DMEM[0] , r_DMEM_ack, 
        \r_WB[4] , \r_WB[3] , \r_WB[2] , \r_WB[1] , \r_WB[0] , r_WB_ack, 
        real_r_WB_ack, real_r_DMEM_ack, real_r_IMEM_ack, n1, n2, n3, n4, n5, 
        n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16;
    wire SYNOPSYS_UNCONNECTED_1 , SYNOPSYS_UNCONNECTED_2 , 
	SYNOPSYS_UNCONNECTED_3 , SYNOPSYS_UNCONNECTED_4 , SYNOPSYS_UNCONNECTED_5 , 
	SYNOPSYS_UNCONNECTED_6 , SYNOPSYS_UNCONNECTED_7 , SYNOPSYS_UNCONNECTED_8 , 
	SYNOPSYS_UNCONNECTED_9 , SYNOPSYS_UNCONNECTED_10 , SYNOPSYS_UNCONNECTED_11 , 
	SYNOPSYS_UNCONNECTED_12 , SYNOPSYS_UNCONNECTED_13 , SYNOPSYS_UNCONNECTED_14 , 
	SYNOPSYS_UNCONNECTED_15 , SYNOPSYS_UNCONNECTED_16 , SYNOPSYS_UNCONNECTED_17 , 
	SYNOPSYS_UNCONNECTED_18 , SYNOPSYS_UNCONNECTED_19 , SYNOPSYS_UNCONNECTED_20 ;
    assign ip_r_sel[3] = 1'b0;
    assign ip_r_sel[2] = 1'b0;
    assign ip_r_sel[1] = 1'b0;
    assign ip_r_sel[0] = 1'b0;
    assign dp_r_sel[3] = 1'b0;
    assign dp_r_sel[2] = 1'b0;
    assign dp_r_sel[1] = 1'b0;
    assign dp_r_sel[0] = 1'b0;
    master_if_iport iport ( .nReset(n1), .mc_req(ip_c_req), .mc_we(ip_c_we), 
        .mc_mult(ip_c_mult), .mc_prd(ip_c_prd), .mc_seq(ip_c_seq), .mc_ts(
        ip_c_ts), .mc_sel(ip_c_sel), .mc_adr(ip_c_adr), .mc_dat(ip_c_dat), 
        .mc_ack(ip_c_ack), .mr_req(ip_r_req), .mr_we(ip_r_we), .mr_err(
        ip_r_err), .mr_rty(ip_r_rty), .mr_acc(ip_r_acc), .mr_ts(ip_r_ts), 
        .mr_dat(ip_r_dat), .mr_ack(ip_r_ack), .chaincommand({\c_Iport[4] , 
        \c_Iport[3] , \c_Iport[2] , \c_Iport[1] , \c_Iport[0] }), 
        .nchaincommandack(real_c_Iport_ack), .chainresponse({\r_Iport[4] , 
        \r_Iport[3] , \r_Iport[2] , \r_Iport[1] , \r_Iport[0] }), 
        .nchainresponseack(r_Iport_ack), .e_bare({1'b0, 1'b0, 1'b1, 1'b0}), 
        .e_dm({1'b0, 1'b0, 1'b0, 1'b1}), .e_im({1'b0, 1'b0, 1'b0, 1'b1}), 
        .e_wish({1'b0, 1'b1, 1'b0, 1'b0}), .r_bare({1'b1, 1'b0, 1'b0, 1'b0}), 
        .r_dm({1'b1, 1'b1, 1'b1, 1'b0}), .r_im({1'b1, 1'b1, 1'b0, 1'b0}), 
        .r_wish({1'b0, 1'b0, 1'b0, 1'b0}), .tag_id({1'b1, 1'b0, 1'b0, 1'b0, 
        1'b0}), .force_bare(force_bare) );
    master_if_dport dport ( .nReset(n3), .mc_req(dp_c_req), .mc_we(dp_c_we), 
        .mc_mult(dp_c_mult), .mc_prd(dp_c_prd), .mc_seq(dp_c_seq), .mc_ts(
        dp_c_ts), .mc_sel(dp_c_sel), .mc_adr(dp_c_adr), .mc_dat(dp_c_dat), 
        .mc_ack(dp_c_ack), .mr_req(dp_r_req), .mr_we(dp_r_we), .mr_err(
        dp_r_err), .mr_rty(dp_r_rty), .mr_acc(dp_r_acc), .mr_ts(dp_r_ts), 
        .mr_dat(dp_r_dat), .mr_ack(dp_r_ack), .chaincommand({\c_Dport[4] , 
        \c_Dport[3] , \c_Dport[2] , \c_Dport[1] , \c_Dport[0] }), 
        .nchaincommandack(real_c_Dport_ack), .chainresponse({\r_Dport[4] , 
        \r_Dport[3] , \r_Dport[2] , \r_Dport[1] , \r_Dport[0] }), 
        .nchainresponseack(r_Dport_ack), .e_bare({1'b0, 1'b0, 1'b1, 1'b0}), 
        .e_dm({1'b0, 1'b0, 1'b0, 1'b1}), .e_im({1'b0, 1'b0, 1'b0, 1'b1}), 
        .e_wish({1'b0, 1'b1, 1'b0, 1'b0}), .r_bare({1'b1, 1'b0, 1'b0, 1'b0}), 
        .r_dm({1'b1, 1'b1, 1'b1, 1'b0}), .r_im({1'b1, 1'b1, 1'b0, 1'b0}), 
        .r_wish({1'b0, 1'b0, 1'b0, 1'b0}), .tag_id({1'b0, 1'b1, 1'b0, 1'b0, 
        1'b0}), .force_bare(force_bare) );
    master_if_tic tic ( .nReset(n3), .mc_req(tic_c_req), .mc_we(tic_c_we), 
        .mc_mult(1'b0), .mc_prd(1'b0), .mc_seq(1'b0), .mc_ts({1'b0, 1'b0, 1'b0
        }), .mc_sel({1'b1, 1'b1, 1'b1, 1'b1}), .mc_adr({\tic_c_adr[31] , 
        \tic_c_adr[30] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \tic_c_adr[11] , 
        \tic_c_adr[10] , \tic_c_adr[9] , \tic_c_adr[8] , \tic_c_adr[7] , 
        \tic_c_adr[6] , \tic_c_adr[5] , \tic_c_adr[4] , \tic_c_adr[3] , 
        \tic_c_adr[2] , 1'b0, 1'b0}), .mc_dat({\tic_c_dat[31] , 
        \tic_c_dat[30] , \tic_c_dat[29] , \tic_c_dat[28] , \tic_c_dat[27] , 
        \tic_c_dat[26] , \tic_c_dat[25] , \tic_c_dat[24] , \tic_c_dat[23] , 
        \tic_c_dat[22] , \tic_c_dat[21] , \tic_c_dat[20] , \tic_c_dat[19] , 
        \tic_c_dat[18] , \tic_c_dat[17] , \tic_c_dat[16] , \tic_c_dat[15] , 
        \tic_c_dat[14] , \tic_c_dat[13] , \tic_c_dat[12] , \tic_c_dat[11] , 
        \tic_c_dat[10] , \tic_c_dat[9] , \tic_c_dat[8] , \tic_c_dat[7] , 
        \tic_c_dat[6] , \tic_c_dat[5] , \tic_c_dat[4] , \tic_c_dat[3] , 
        \tic_c_dat[2] , \tic_c_dat[1] , \tic_c_dat[0] }), .mc_ack(tic_c_ack), 
        .mr_req(tic_r_req), .mr_dat({\tic_r_dat[31] , \tic_r_dat[30] , 
        \tic_r_dat[29] , \tic_r_dat[28] , \tic_r_dat[27] , \tic_r_dat[26] , 
        \tic_r_dat[25] , \tic_r_dat[24] , \tic_r_dat[23] , \tic_r_dat[22] , 
        \tic_r_dat[21] , \tic_r_dat[20] , \tic_r_dat[19] , \tic_r_dat[18] , 
        \tic_r_dat[17] , \tic_r_dat[16] , \tic_r_dat[15] , \tic_r_dat[14] , 
        \tic_r_dat[13] , \tic_r_dat[12] , \tic_r_dat[11] , \tic_r_dat[10] , 
        \tic_r_dat[9] , \tic_r_dat[8] , \tic_r_dat[7] , \tic_r_dat[6] , 
        \tic_r_dat[5] , \tic_r_dat[4] , \tic_r_dat[3] , \tic_r_dat[2] , 
        \tic_r_dat[1] , \tic_r_dat[0] }), .mr_ack(tic_r_ack), .chaincommand({
        \c_TIC[4] , \c_TIC[3] , \c_TIC[2] , \c_TIC[1] , \c_TIC[0] }), 
        .nchaincommandack(real_c_TIC_ack), .chainresponse({\r_TIC[4] , 
        \r_TIC[3] , \r_TIC[2] , \r_TIC[1] , \r_TIC[0] }), .nchainresponseack(
        r_TIC_ack), .e_bare({1'b0, 1'b0, 1'b1, 1'b0}), .e_dm({1'b0, 1'b0, 1'b0, 
        1'b1}), .e_im({1'b0, 1'b0, 1'b0, 1'b1}), .e_wish({1'b0, 1'b1, 1'b0, 
        1'b0}), .r_bare({1'b1, 1'b0, 1'b0, 1'b0}), .r_dm({1'b1, 1'b1, 1'b1, 
        1'b0}), .r_im({1'b1, 1'b1, 1'b0, 1'b0}), .r_wish({1'b0, 1'b0, 1'b0, 
        1'b0}), .tag_id({1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .force_bare(
        force_bare) );
    tic ticBlock ( .c_req(ei_c_req), .c_ack(ei_c_ack), .c_we(ei_c_we), 
        .c_addr(ei_c_addr), .r_req(ei_r_req), .r_ack(ei_r_ack), .data_in(
        ei_data_in), .data_out(ei_data_out), .reset_b(n4), .mc_req(tic_c_req), 
        .mc_we(tic_c_we), .mc_adr({\tic_c_adr[31] , \tic_c_adr[30] , 
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, \tic_c_adr[11] , \tic_c_adr[10] , 
        \tic_c_adr[9] , \tic_c_adr[8] , \tic_c_adr[7] , \tic_c_adr[6] , 
        \tic_c_adr[5] , \tic_c_adr[4] , \tic_c_adr[3] , \tic_c_adr[2] , 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20}), .mc_dat({
        \tic_c_dat[31] , \tic_c_dat[30] , \tic_c_dat[29] , \tic_c_dat[28] , 
        \tic_c_dat[27] , \tic_c_dat[26] , \tic_c_dat[25] , \tic_c_dat[24] , 
        \tic_c_dat[23] , \tic_c_dat[22] , \tic_c_dat[21] , \tic_c_dat[20] , 
        \tic_c_dat[19] , \tic_c_dat[18] , \tic_c_dat[17] , \tic_c_dat[16] , 
        \tic_c_dat[15] , \tic_c_dat[14] , \tic_c_dat[13] , \tic_c_dat[12] , 
        \tic_c_dat[11] , \tic_c_dat[10] , \tic_c_dat[9] , \tic_c_dat[8] , 
        \tic_c_dat[7] , \tic_c_dat[6] , \tic_c_dat[5] , \tic_c_dat[4] , 
        \tic_c_dat[3] , \tic_c_dat[2] , \tic_c_dat[1] , \tic_c_dat[0] }), 
        .mc_ack(tic_c_ack), .mr_req(tic_r_req), .mr_dat({\tic_r_dat[31] , 
        \tic_r_dat[30] , \tic_r_dat[29] , \tic_r_dat[28] , \tic_r_dat[27] , 
        \tic_r_dat[26] , \tic_r_dat[25] , \tic_r_dat[24] , \tic_r_dat[23] , 
        \tic_r_dat[22] , \tic_r_dat[21] , \tic_r_dat[20] , \tic_r_dat[19] , 
        \tic_r_dat[18] , \tic_r_dat[17] , \tic_r_dat[16] , \tic_r_dat[15] , 
        \tic_r_dat[14] , \tic_r_dat[13] , \tic_r_dat[12] , \tic_r_dat[11] , 
        \tic_r_dat[10] , \tic_r_dat[9] , \tic_r_dat[8] , \tic_r_dat[7] , 
        \tic_r_dat[6] , \tic_r_dat[5] , \tic_r_dat[4] , \tic_r_dat[3] , 
        \tic_r_dat[2] , \tic_r_dat[1] , \tic_r_dat[0] }), .mr_ack(tic_r_ack)
         );
    inv_2 U10 ( .x(c_BC_ack_n), .a(c_BC_ack) );
    inv_2 U12 ( .x(c_WB_ack_n), .a(c_WB_ack) );
    inv_2 U13 ( .x(c_IMEM_ack_n), .a(c_IMEM_ack) );
    inv_2 U14 ( .x(c_DMEM_ack_n), .a(c_DMEM_ack) );
    comm_fab_scan cmd_fab ( .nrst(n2), .I_port_eop_i(\c_Iport[4] ), 
        .I_port_d0_i(\c_Iport[0] ), .I_port_d1_i(\c_Iport[1] ), .I_port_d2_i(
        \c_Iport[2] ), .I_port_d3_i(\c_Iport[3] ), .I_port_ack(c_Iport_ack), 
        .TIC_eop_i(\c_TIC[4] ), .TIC_d0_i(\c_TIC[0] ), .TIC_d1_i(\c_TIC[1] ), 
        .TIC_d2_i(\c_TIC[2] ), .TIC_d3_i(\c_TIC[3] ), .TIC_ack(c_TIC_ack), 
        .D_port_eop_i(\c_Dport[4] ), .D_port_d0_i(\c_Dport[0] ), .D_port_d1_i(
        \c_Dport[1] ), .D_port_d2_i(\c_Dport[2] ), .D_port_d3_i(\c_Dport[3] ), 
        .D_port_ack(c_Dport_ack), .BC_eop_i(c_BC[4]), .BC_d0_i(c_BC[0]), 
        .BC_d1_i(c_BC[1]), .BC_d2_i(c_BC[2]), .BC_d3_i(c_BC[3]), .BC_ack(
        c_BC_ack_n), .WB_eop_i(\c_WB[4] ), .WB_d0_i(\c_WB[0] ), .WB_d1_i(
        \c_WB[1] ), .WB_d2_i(\c_WB[2] ), .WB_d3_i(\c_WB[3] ), .WB_ack(
        c_WB_ack_n), .IMEM_eop_i(\c_IMEM[4] ), .IMEM_d0_i(\c_IMEM[0] ), 
        .IMEM_d1_i(\c_IMEM[1] ), .IMEM_d2_i(\c_IMEM[2] ), .IMEM_d3_i(
        \c_IMEM[3] ), .IMEM_ack(c_IMEM_ack_n), .DMEM_eop_i(\c_DMEM[4] ), 
        .DMEM_d0_i(\c_DMEM[0] ), .DMEM_d1_i(\c_DMEM[1] ), .DMEM_d2_i(
        \c_DMEM[2] ), .DMEM_d3_i(\c_DMEM[3] ), .DMEM_ack(c_DMEM_ack_n), 
        .test_si(test_si), .test_so(scan_o_cmd), .test_se(n12), .phi1(n9), 
        .phi2(n15), .phi3(n6) );
    inv_2 U20 ( .x(r_Iport_ack_n), .a(r_Iport_ack) );
    inv_2 U21 ( .x(r_TIC_ack_n), .a(r_TIC_ack) );
    inv_2 U22 ( .x(r_Dport_ack_n), .a(r_Dport_ack) );
    resp_fab_scan rsp_fab ( .nrst(n3), .IMEM_eop_i(\r_IMEM[4] ), .IMEM_d0_i(
        \r_IMEM[0] ), .IMEM_d1_i(\r_IMEM[1] ), .IMEM_d2_i(\r_IMEM[2] ), 
        .IMEM_d3_i(\r_IMEM[3] ), .IMEM_ack(r_IMEM_ack), .DMEM_eop_i(
        \r_DMEM[4] ), .DMEM_d0_i(\r_DMEM[0] ), .DMEM_d1_i(\r_DMEM[1] ), 
        .DMEM_d2_i(\r_DMEM[2] ), .DMEM_d3_i(\r_DMEM[3] ), .DMEM_ack(r_DMEM_ack
        ), .WB_eop_i(\r_WB[4] ), .WB_d0_i(\r_WB[0] ), .WB_d1_i(\r_WB[1] ), 
        .WB_d2_i(\r_WB[2] ), .WB_d3_i(\r_WB[3] ), .WB_ack(r_WB_ack), 
        .BC_eop_i(r_BC[4]), .BC_d0_i(r_BC[0]), .BC_d1_i(r_BC[1]), .BC_d2_i(
        r_BC[2]), .BC_d3_i(r_BC[3]), .BC_ack(r_BC_ack), .I_port_eop_i(
        \r_Iport[4] ), .I_port_d0_i(\r_Iport[0] ), .I_port_d1_i(\r_Iport[1] ), 
        .I_port_d2_i(\r_Iport[2] ), .I_port_d3_i(\r_Iport[3] ), .I_port_ack(
        r_Iport_ack_n), .TIC_eop_i(\r_TIC[4] ), .TIC_d0_i(\r_TIC[0] ), 
        .TIC_d1_i(\r_TIC[1] ), .TIC_d2_i(\r_TIC[2] ), .TIC_d3_i(\r_TIC[3] ), 
        .TIC_ack(r_TIC_ack_n), .D_port_eop_i(\r_Dport[4] ), .D_port_d0_i(
        \r_Dport[0] ), .D_port_d1_i(\r_Dport[1] ), .D_port_d2_i(\r_Dport[2] ), 
        .D_port_d3_i(\r_Dport[3] ), .D_port_ack(r_Dport_ack_n), .test_si(
        scan_o_cmd), .test_so(test_so), .test_se(n13), .phi1(n10), .phi2(n16), 
        .phi3(n7) );
    wb_block wb ( .nReset(n1), .clk(clk), .chaincommand({\c_WB[4] , \c_WB[3] , 
        \c_WB[2] , \c_WB[1] , \c_WB[0] }), .nchaincommandack(c_WB_ack), 
        .chainresponse({\r_WB[4] , \r_WB[3] , \r_WB[2] , \r_WB[1] , \r_WB[0] }
        ), .nchainresponseack(real_r_WB_ack), .e_dp({1'b0, 1'b0, 1'b1}), 
        .e_ip({1'b0, 1'b0, 1'b1}), .e_tic({1'b0, 1'b1, 1'b0}), .r_dp({1'b1, 
        1'b0, 1'b0}), .r_ip({1'b1, 1'b1, 1'b0}), .r_tic({1'b0, 1'b0, 1'b0}), 
        .wb_we_o(wish_we_o), .wb_stb_cyc_o(wish_stb_cyc_o), .wb_ack_i(
        wish_ack_i), .wb_adr_o(wish_adr_o), .wb_dat_i(wish_dat_i), .wb_dat_o(
        wish_dat_o) );
    slave_if_dmem dmem ( .nReset(n1), .sc_req(dm_c_req), .sc_we(dm_c_we), 
        .sc_mult(dm_c_mult), .sc_seq(dm_c_seq), .sc_prd(dm_c_prd), .sc_ts(
        dm_c_ts), .sc_st(dm_c_st), .sc_sel(dm_c_sel), .sc_adr(dm_c_adr), 
        .sc_dat(dm_c_dat), .sc_ack(dm_c_ack), .sr_req(dm_r_req), .sr_err(
        dm_r_err), .sr_rty(dm_r_rty), .sr_acc(dm_r_acc), .sr_mult(dm_r_mult), 
        .sr_ts(dm_r_ts), .sr_rt(dm_r_rt), .sr_sel(dm_r_sel), .sr_dat(dm_r_dat), 
        .sr_ack(dm_r_ack), .chaincommand({\c_DMEM[4] , \c_DMEM[3] , 
        \c_DMEM[2] , \c_DMEM[1] , \c_DMEM[0] }), .nchaincommandack(c_DMEM_ack), 
        .chainresponse({\r_DMEM[4] , \r_DMEM[3] , \r_DMEM[2] , \r_DMEM[1] , 
        \r_DMEM[0] }), .nchainresponseack(real_r_DMEM_ack), .e_dp({1'b0, 1'b0, 
        1'b1}), .e_ip({1'b0, 1'b0, 1'b1}), .e_tic({1'b0, 1'b1, 1'b0}), .r_dp({
        1'b1, 1'b0, 1'b0}), .r_ip({1'b1, 1'b1, 1'b0}), .r_tic({1'b0, 1'b0, 
        1'b0}) );
    slave_if_imem imem ( .nReset(n4), .sc_req(im_c_req), .sc_we(im_c_we), 
        .sc_mult(im_c_mult), .sc_seq(im_c_seq), .sc_prd(im_c_prd), .sc_ts(
        im_c_ts), .sc_st(im_c_st), .sc_sel(im_c_sel), .sc_adr(im_c_adr), 
        .sc_dat(im_c_dat), .sc_ack(im_c_ack), .sr_req(im_r_req), .sr_err(
        im_r_err), .sr_rty(im_r_rty), .sr_acc(im_r_acc), .sr_mult(im_r_mult), 
        .sr_ts(im_r_ts), .sr_rt(im_r_rt), .sr_sel(im_r_sel), .sr_dat(im_r_dat), 
        .sr_ack(im_r_ack), .chaincommand({\c_IMEM[4] , \c_IMEM[3] , 
        \c_IMEM[2] , \c_IMEM[1] , \c_IMEM[0] }), .nchaincommandack(c_IMEM_ack), 
        .chainresponse({\r_IMEM[4] , \r_IMEM[3] , \r_IMEM[2] , \r_IMEM[1] , 
        \r_IMEM[0] }), .nchainresponseack(real_r_IMEM_ack), .e_dp({1'b0, 1'b0, 
        1'b1}), .e_ip({1'b0, 1'b0, 1'b1}), .e_tic({1'b0, 1'b1, 1'b0}), .r_dp({
        1'b1, 1'b0, 1'b0}), .r_ip({1'b1, 1'b1, 1'b0}), .r_tic({1'b0, 1'b0, 
        1'b0}) );
    inv_2 U8 ( .x(n6), .a(n5) );
    inv_2 U9 ( .x(n7), .a(n5) );
    inv_2 U11 ( .x(n15), .a(n14) );
    inv_2 U15 ( .x(n13), .a(n11) );
    inv_2 U16 ( .x(n9), .a(n8) );
    inv_2 U17 ( .x(n10), .a(n8) );
    inv_2 U18 ( .x(n12), .a(n11) );
    inv_2 U19 ( .x(n16), .a(n14) );
    buf_3 U23 ( .x(n1), .a(nrst) );
    buf_3 U24 ( .x(n4), .a(nrst) );
    buf_4 U25 ( .x(n2), .a(nrst) );
    buf_4 U26 ( .x(n3), .a(nrst) );
    inv_2 U27 ( .x(n5), .a(phi3) );
    inv_2 U28 ( .x(n8), .a(phi1) );
    inv_5 U29 ( .x(n11), .a(test_se) );
    inv_2 U30 ( .x(n14), .a(phi2) );
    inv_5 U31 ( .x(rst), .a(n4) );
    nor2_4 U32 ( .x(real_c_Dport_ack), .a(rst), .b(c_Dport_ack) );
    nor2_4 U33 ( .x(real_r_IMEM_ack), .a(rst), .b(r_IMEM_ack) );
    nor2_4 U34 ( .x(real_r_DMEM_ack), .a(rst), .b(r_DMEM_ack) );
    nor2_4 U35 ( .x(real_r_WB_ack), .a(rst), .b(r_WB_ack) );
    nor2_4 U36 ( .x(real_c_TIC_ack), .a(rst), .b(c_TIC_ack) );
    nor2_4 U37 ( .x(real_c_Iport_ack), .a(rst), .b(c_Iport_ack) );
endmodule


module aspida_net ( nrst_pad, clk_pad, ip_c_req, ip_c_we, ip_c_mult, ip_c_prd, 
    ip_c_seq, ip_c_ts, ip_c_sel, ip_c_adr, ip_c_dat, ip_c_ack, ip_r_req, 
    ip_r_we, ip_r_err, ip_r_rty, ip_r_acc, ip_r_ts, ip_r_sel, ip_r_dat, 
    ip_r_ack, dp_c_req, dp_c_we, dp_c_mult, dp_c_prd, dp_c_seq, dp_c_ts, 
    dp_c_sel, dp_c_adr, dp_c_dat, dp_c_ack, dp_r_req, dp_r_we, dp_r_err, 
    dp_r_rty, dp_r_acc, dp_r_ts, dp_r_sel, dp_r_dat, dp_r_ack, ei_c_req_pad, 
    ei_c_ack_pad, ei_c_we_pad, ei_c_addr_pad, ei_r_req_pad, ei_r_ack_pad, 
    ei_data_pad, c_BC_pad, c_BC_ack_pad, r_BC_pad, r_BC_ack_pad, wish_we_o_pad, 
    wish_stb_cyc_o_pad, wish_ack_i_pad, wish_adr_o_pad, wish_dat_pad, dm_c_req, 
    dm_c_we, dm_c_mult, dm_c_seq, dm_c_prd, dm_c_ts, dm_c_st, dm_c_sel, 
    dm_c_adr, dm_c_dat, dm_c_ack, dm_r_req, dm_r_err, dm_r_rty, dm_r_acc, 
    dm_r_mult, dm_r_ts, dm_r_rt, dm_r_sel, dm_r_dat, dm_r_ack, im_c_req, 
    im_c_we, im_c_mult, im_c_seq, im_c_prd, im_c_ts, im_c_st, im_c_sel, 
    im_c_adr, im_c_dat, im_c_ack, im_r_req, im_r_err, im_r_rty, im_r_acc, 
    im_r_mult, im_r_ts, im_r_rt, im_r_sel, im_r_dat, im_r_ack, test_si_pad, 
    test_so_pad, test_se_pad, phi1_pad, phi2_pad, phi3_pad, force_bare_pad );
input  [2:0] ip_c_ts;
input  [3:0] ip_c_sel;
input  [31:0] ip_c_adr;
input  [31:0] ip_c_dat;
output [2:0] ip_r_ts;
output [3:0] ip_r_sel;
output [31:0] ip_r_dat;
input  [2:0] dp_c_ts;
input  [3:0] dp_c_sel;
input  [31:0] dp_c_adr;
input  [31:0] dp_c_dat;
output [2:0] dp_r_ts;
output [3:0] dp_r_sel;
output [31:0] dp_r_dat;
input  [10:0] ei_c_addr_pad;
inout  [7:0] ei_data_pad;
output [4:0] c_BC_pad;
input  [4:0] r_BC_pad;
output [11:0] wish_adr_o_pad;
inout  [31:0] wish_dat_pad;
output [2:0] dm_c_ts;
output [4:0] dm_c_st;
output [3:0] dm_c_sel;
output [31:0] dm_c_adr;
output [31:0] dm_c_dat;
input  [2:0] dm_r_ts;
input  [4:0] dm_r_rt;
input  [3:0] dm_r_sel;
input  [31:0] dm_r_dat;
output [2:0] im_c_ts;
output [4:0] im_c_st;
output [3:0] im_c_sel;
output [31:0] im_c_adr;
output [31:0] im_c_dat;
input  [2:0] im_r_ts;
input  [4:0] im_r_rt;
input  [3:0] im_r_sel;
input  [31:0] im_r_dat;
input  nrst_pad, clk_pad, ip_c_req, ip_c_we, ip_c_mult, ip_c_prd, ip_c_seq, 
    ip_r_ack, dp_c_req, dp_c_we, dp_c_mult, dp_c_prd, dp_c_seq, dp_r_ack, 
    ei_c_req_pad, ei_c_we_pad, ei_r_ack_pad, c_BC_ack_pad, wish_ack_i_pad, 
    dm_c_ack, dm_r_req, dm_r_err, dm_r_rty, dm_r_acc, dm_r_mult, im_c_ack, 
    im_r_req, im_r_err, im_r_rty, im_r_acc, im_r_mult, test_si_pad, 
    test_se_pad, phi1_pad, phi2_pad, phi3_pad, force_bare_pad;
output ip_c_ack, ip_r_req, ip_r_we, ip_r_err, ip_r_rty, ip_r_acc, dp_c_ack, 
    dp_r_req, dp_r_we, dp_r_err, dp_r_rty, dp_r_acc, ei_c_ack_pad, 
    ei_r_req_pad, r_BC_ack_pad, wish_we_o_pad, wish_stb_cyc_o_pad, dm_c_req, 
    dm_c_we, dm_c_mult, dm_c_seq, dm_c_prd, dm_r_ack, im_c_req, im_c_we, 
    im_c_mult, im_c_seq, im_c_prd, im_r_ack, test_so_pad;
    wire nrst, clk, ei_c_req, ei_c_ack, ei_c_we, \ei_c_addr[10] , 
        \ei_c_addr[9] , \ei_c_addr[8] , \ei_c_addr[7] , \ei_c_addr[6] , 
        \ei_c_addr[5] , \ei_c_addr[4] , \ei_c_addr[3] , \ei_c_addr[2] , 
        \ei_c_addr[1] , \ei_c_addr[0] , ei_r_req, ei_r_ack, \c_BC[4] , 
        \c_BC[3] , \c_BC[2] , \c_BC[1] , \c_BC[0] , c_BC_ack, \r_BC[4] , 
        \r_BC[3] , \r_BC[2] , \r_BC[1] , \r_BC[0] , r_BC_ack, wish_we_o, 
        wish_stb_cyc_o, wish_ack_i, \wish_adr_o[11] , \wish_adr_o[10] , 
        \wish_adr_o[9] , \wish_adr_o[8] , \wish_adr_o[7] , \wish_adr_o[6] , 
        \wish_adr_o[5] , \wish_adr_o[4] , \wish_adr_o[3] , \wish_adr_o[2] , 
        \wish_adr_o[1] , \wish_adr_o[0] , test_si, test_se, phi1, phi2, phi3, 
        test_so, force_bare, \ei_data_in[7] , \ei_data_in[6] , \ei_data_in[5] , 
        \ei_data_in[4] , \ei_data_in[3] , \ei_data_in[2] , \ei_data_in[1] , 
        \ei_data_in[0] , \ei_data_out[7] , \ei_data_out[6] , \ei_data_out[5] , 
        \ei_data_out[4] , \ei_data_out[3] , \ei_data_out[2] , \ei_data_out[1] , 
        \ei_data_out[0] , \wish_dat_i[31] , \wish_dat_i[30] , \wish_dat_i[29] , 
        \wish_dat_i[28] , \wish_dat_i[27] , \wish_dat_i[26] , \wish_dat_i[25] , 
        \wish_dat_i[24] , \wish_dat_i[23] , \wish_dat_i[22] , \wish_dat_i[21] , 
        \wish_dat_i[20] , \wish_dat_i[19] , \wish_dat_i[18] , \wish_dat_i[17] , 
        \wish_dat_i[16] , \wish_dat_i[15] , \wish_dat_i[14] , \wish_dat_i[13] , 
        \wish_dat_i[12] , \wish_dat_i[11] , \wish_dat_i[10] , \wish_dat_i[9] , 
        \wish_dat_i[8] , \wish_dat_i[7] , \wish_dat_i[6] , \wish_dat_i[5] , 
        \wish_dat_i[4] , \wish_dat_i[3] , \wish_dat_i[2] , \wish_dat_i[1] , 
        \wish_dat_i[0] , \wish_dat_o[31] , \wish_dat_o[30] , \wish_dat_o[29] , 
        \wish_dat_o[28] , \wish_dat_o[27] , \wish_dat_o[26] , \wish_dat_o[25] , 
        \wish_dat_o[24] , \wish_dat_o[23] , \wish_dat_o[22] , \wish_dat_o[21] , 
        \wish_dat_o[20] , \wish_dat_o[19] , \wish_dat_o[18] , \wish_dat_o[17] , 
        \wish_dat_o[16] , \wish_dat_o[15] , \wish_dat_o[14] , \wish_dat_o[13] , 
        \wish_dat_o[12] , \wish_dat_o[11] , \wish_dat_o[10] , \wish_dat_o[9] , 
        \wish_dat_o[8] , \wish_dat_o[7] , \wish_dat_o[6] , \wish_dat_o[5] , 
        \wish_dat_o[4] , \wish_dat_o[3] , \wish_dat_o[2] , \wish_dat_o[1] , 
        \wish_dat_o[0] , ei_c_we_b;
    inbuf3_16 reset_pad ( .di(nrst), .pad(nrst_pad) );
    inv_4 U3 ( .x(ei_c_we_b), .a(ei_c_we) );
    inbuf3_16 ticCreq_pad ( .di(ei_c_req), .pad(ei_c_req_pad) );
    iobuf2_16_4 ticCack_pad ( .pad(ei_c_ack_pad), .\do (ei_c_ack), .en(1'b1)
         );
    inbuf3_16 ticWe_pad ( .di(ei_c_we), .pad(ei_c_we_pad) );
    inbuf3_16 ticAddr_0_pad ( .di(\ei_c_addr[0] ), .pad(ei_c_addr_pad[0]) );
    inbuf3_16 ticAddr_1_pad ( .di(\ei_c_addr[1] ), .pad(ei_c_addr_pad[1]) );
    inbuf3_16 ticAddr_2_pad ( .di(\ei_c_addr[2] ), .pad(ei_c_addr_pad[2]) );
    inbuf3_16 ticAddr_3_pad ( .di(\ei_c_addr[3] ), .pad(ei_c_addr_pad[3]) );
    inbuf3_16 ticAddr_4_pad ( .di(\ei_c_addr[4] ), .pad(ei_c_addr_pad[4]) );
    inbuf3_16 ticAddr_5_pad ( .di(\ei_c_addr[5] ), .pad(ei_c_addr_pad[5]) );
    inbuf3_16 ticAddr_6_pad ( .di(\ei_c_addr[6] ), .pad(ei_c_addr_pad[6]) );
    inbuf3_16 ticAddr_7_pad ( .di(\ei_c_addr[7] ), .pad(ei_c_addr_pad[7]) );
    inbuf3_16 ticAddr_8_pad ( .di(\ei_c_addr[8] ), .pad(ei_c_addr_pad[8]) );
    inbuf3_16 ticAddr_9_pad ( .di(\ei_c_addr[9] ), .pad(ei_c_addr_pad[9]) );
    inbuf3_16 ticAddr_10_pad ( .di(\ei_c_addr[10] ), .pad(ei_c_addr_pad[10])
         );
    iobuf2_16_4 ticRreq_pad ( .pad(ei_r_req_pad), .\do (ei_r_req), .en(1'b1)
         );
    inbuf3_16 ticRack_pad ( .di(ei_r_ack), .pad(ei_r_ack_pad) );
    iobuf3_16_4 tic_dat_pad_0 ( .di(\ei_data_in[0] ), .pad(ei_data_pad[0]), 
        .\do (\ei_data_out[0] ), .en(ei_c_we_b) );
    iobuf3_16_4 tic_dat_pad_1 ( .di(\ei_data_in[1] ), .pad(ei_data_pad[1]), 
        .\do (\ei_data_out[1] ), .en(ei_c_we_b) );
    iobuf3_16_4 tic_dat_pad_2 ( .di(\ei_data_in[2] ), .pad(ei_data_pad[2]), 
        .\do (\ei_data_out[2] ), .en(ei_c_we_b) );
    iobuf3_16_4 tic_dat_pad_3 ( .di(\ei_data_in[3] ), .pad(ei_data_pad[3]), 
        .\do (\ei_data_out[3] ), .en(ei_c_we_b) );
    iobuf3_16_4 tic_dat_pad_4 ( .di(\ei_data_in[4] ), .pad(ei_data_pad[4]), 
        .\do (\ei_data_out[4] ), .en(ei_c_we_b) );
    iobuf3_16_4 tic_dat_pad_5 ( .di(\ei_data_in[5] ), .pad(ei_data_pad[5]), 
        .\do (\ei_data_out[5] ), .en(ei_c_we_b) );
    iobuf3_16_4 tic_dat_pad_6 ( .di(\ei_data_in[6] ), .pad(ei_data_pad[6]), 
        .\do (\ei_data_out[6] ), .en(ei_c_we_b) );
    iobuf3_16_4 tic_dat_pad_7 ( .di(\ei_data_in[7] ), .pad(ei_data_pad[7]), 
        .\do (\ei_data_out[7] ), .en(ei_c_we_b) );
    iobuf2_16_4 bc_Cpad_0 ( .pad(c_BC_pad[0]), .\do (\c_BC[0] ), .en(1'b1) );
    iobuf2_16_4 bc_Cpad_1 ( .pad(c_BC_pad[1]), .\do (\c_BC[1] ), .en(1'b1) );
    iobuf2_16_4 bc_Cpad_2 ( .pad(c_BC_pad[2]), .\do (\c_BC[2] ), .en(1'b1) );
    iobuf2_16_4 bc_Cpad_3 ( .pad(c_BC_pad[3]), .\do (\c_BC[3] ), .en(1'b1) );
    iobuf2_16_4 bc_Cpad_4 ( .pad(c_BC_pad[4]), .\do (\c_BC[4] ), .en(1'b1) );
    inbuf3_16 bc_Cack_pad ( .di(c_BC_ack), .pad(c_BC_ack_pad) );
    inbuf3_16 bc_Rpad_0 ( .di(\r_BC[0] ), .pad(r_BC_pad[0]) );
    inbuf3_16 bc_Rpad_1 ( .di(\r_BC[1] ), .pad(r_BC_pad[1]) );
    inbuf3_16 bc_Rpad_2 ( .di(\r_BC[2] ), .pad(r_BC_pad[2]) );
    inbuf3_16 bc_Rpad_3 ( .di(\r_BC[3] ), .pad(r_BC_pad[3]) );
    inbuf3_16 bc_Rpad_4 ( .di(\r_BC[4] ), .pad(r_BC_pad[4]) );
    iobuf2_16_4 bc_Rack_pad ( .pad(r_BC_ack_pad), .\do (r_BC_ack), .en(1'b1)
         );
    inbuf3_16 clock_pad ( .di(clk), .pad(clk_pad) );
    iobuf2_16_4 wb_we_pad ( .pad(wish_we_o_pad), .\do (wish_we_o), .en(1'b1)
         );
    iobuf2_16_4 wb_stb_cyc_pad ( .pad(wish_stb_cyc_o_pad), .\do (
        wish_stb_cyc_o), .en(1'b1) );
    inbuf3_16 wb_ack_pad ( .di(wish_ack_i), .pad(wish_ack_i_pad) );
    iobuf2_16_4 wb_adr_pad_0 ( .pad(wish_adr_o_pad[0]), .\do (\wish_adr_o[0] ), 
        .en(1'b1) );
    iobuf2_16_4 wb_adr_pad_1 ( .pad(wish_adr_o_pad[1]), .\do (\wish_adr_o[1] ), 
        .en(1'b1) );
    iobuf2_16_4 wb_adr_pad_2 ( .pad(wish_adr_o_pad[2]), .\do (\wish_adr_o[2] ), 
        .en(1'b1) );
    iobuf2_16_4 wb_adr_pad_3 ( .pad(wish_adr_o_pad[3]), .\do (\wish_adr_o[3] ), 
        .en(1'b1) );
    iobuf2_16_4 wb_adr_pad_4 ( .pad(wish_adr_o_pad[4]), .\do (\wish_adr_o[4] ), 
        .en(1'b1) );
    iobuf2_16_4 wb_adr_pad_5 ( .pad(wish_adr_o_pad[5]), .\do (\wish_adr_o[5] ), 
        .en(1'b1) );
    iobuf2_16_4 wb_adr_pad_6 ( .pad(wish_adr_o_pad[6]), .\do (\wish_adr_o[6] ), 
        .en(1'b1) );
    iobuf2_16_4 wb_adr_pad_7 ( .pad(wish_adr_o_pad[7]), .\do (\wish_adr_o[7] ), 
        .en(1'b1) );
    iobuf2_16_4 wb_adr_pad_8 ( .pad(wish_adr_o_pad[8]), .\do (\wish_adr_o[8] ), 
        .en(1'b1) );
    iobuf2_16_4 wb_adr_pad_9 ( .pad(wish_adr_o_pad[9]), .\do (\wish_adr_o[9] ), 
        .en(1'b1) );
    iobuf2_16_4 wb_adr_pad_10 ( .pad(wish_adr_o_pad[10]), .\do (
        \wish_adr_o[10] ), .en(1'b1) );
    iobuf2_16_4 wb_adr_pad_11 ( .pad(wish_adr_o_pad[11]), .\do (
        \wish_adr_o[11] ), .en(1'b1) );
    iobuf3_16_4 wb_dat_pad_0 ( .di(\wish_dat_i[0] ), .pad(wish_dat_pad[0]), 
        .\do (\wish_dat_o[0] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_1 ( .di(\wish_dat_i[1] ), .pad(wish_dat_pad[1]), 
        .\do (\wish_dat_o[1] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_2 ( .di(\wish_dat_i[2] ), .pad(wish_dat_pad[2]), 
        .\do (\wish_dat_o[2] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_3 ( .di(\wish_dat_i[3] ), .pad(wish_dat_pad[3]), 
        .\do (\wish_dat_o[3] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_4 ( .di(\wish_dat_i[4] ), .pad(wish_dat_pad[4]), 
        .\do (\wish_dat_o[4] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_5 ( .di(\wish_dat_i[5] ), .pad(wish_dat_pad[5]), 
        .\do (\wish_dat_o[5] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_6 ( .di(\wish_dat_i[6] ), .pad(wish_dat_pad[6]), 
        .\do (\wish_dat_o[6] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_7 ( .di(\wish_dat_i[7] ), .pad(wish_dat_pad[7]), 
        .\do (\wish_dat_o[7] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_8 ( .di(\wish_dat_i[8] ), .pad(wish_dat_pad[8]), 
        .\do (\wish_dat_o[8] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_9 ( .di(\wish_dat_i[9] ), .pad(wish_dat_pad[9]), 
        .\do (\wish_dat_o[9] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_10 ( .di(\wish_dat_i[10] ), .pad(wish_dat_pad[10]), 
        .\do (\wish_dat_o[10] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_11 ( .di(\wish_dat_i[11] ), .pad(wish_dat_pad[11]), 
        .\do (\wish_dat_o[11] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_12 ( .di(\wish_dat_i[12] ), .pad(wish_dat_pad[12]), 
        .\do (\wish_dat_o[12] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_13 ( .di(\wish_dat_i[13] ), .pad(wish_dat_pad[13]), 
        .\do (\wish_dat_o[13] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_14 ( .di(\wish_dat_i[14] ), .pad(wish_dat_pad[14]), 
        .\do (\wish_dat_o[14] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_15 ( .di(\wish_dat_i[15] ), .pad(wish_dat_pad[15]), 
        .\do (\wish_dat_o[15] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_16 ( .di(\wish_dat_i[16] ), .pad(wish_dat_pad[16]), 
        .\do (\wish_dat_o[16] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_17 ( .di(\wish_dat_i[17] ), .pad(wish_dat_pad[17]), 
        .\do (\wish_dat_o[17] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_18 ( .di(\wish_dat_i[18] ), .pad(wish_dat_pad[18]), 
        .\do (\wish_dat_o[18] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_19 ( .di(\wish_dat_i[19] ), .pad(wish_dat_pad[19]), 
        .\do (\wish_dat_o[19] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_20 ( .di(\wish_dat_i[20] ), .pad(wish_dat_pad[20]), 
        .\do (\wish_dat_o[20] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_21 ( .di(\wish_dat_i[21] ), .pad(wish_dat_pad[21]), 
        .\do (\wish_dat_o[21] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_22 ( .di(\wish_dat_i[22] ), .pad(wish_dat_pad[22]), 
        .\do (\wish_dat_o[22] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_23 ( .di(\wish_dat_i[23] ), .pad(wish_dat_pad[23]), 
        .\do (\wish_dat_o[23] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_24 ( .di(\wish_dat_i[24] ), .pad(wish_dat_pad[24]), 
        .\do (\wish_dat_o[24] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_25 ( .di(\wish_dat_i[25] ), .pad(wish_dat_pad[25]), 
        .\do (\wish_dat_o[25] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_26 ( .di(\wish_dat_i[26] ), .pad(wish_dat_pad[26]), 
        .\do (\wish_dat_o[26] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_27 ( .di(\wish_dat_i[27] ), .pad(wish_dat_pad[27]), 
        .\do (\wish_dat_o[27] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_28 ( .di(\wish_dat_i[28] ), .pad(wish_dat_pad[28]), 
        .\do (\wish_dat_o[28] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_29 ( .di(\wish_dat_i[29] ), .pad(wish_dat_pad[29]), 
        .\do (\wish_dat_o[29] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_30 ( .di(\wish_dat_i[30] ), .pad(wish_dat_pad[30]), 
        .\do (\wish_dat_o[30] ), .en(wish_we_o) );
    iobuf3_16_4 wb_dat_pad_31 ( .di(\wish_dat_i[31] ), .pad(wish_dat_pad[31]), 
        .\do (\wish_dat_o[31] ), .en(wish_we_o) );
    inbuf3_16 si_pad ( .di(test_si), .pad(test_si_pad) );
    inbuf3_16 se_pad ( .di(test_se), .pad(test_se_pad) );
    inbuf3_16 phi_1_pad ( .di(phi1), .pad(phi1_pad) );
    inbuf3_16 phi_2_pad ( .di(phi2), .pad(phi2_pad) );
    inbuf3_16 phi_3_pad ( .di(phi3), .pad(phi3_pad) );
    iobuf3_16_4 so_pad ( .pad(test_so_pad), .\do (test_so), .en(1'b1) );
    inbuf3_16 forceBC_pad ( .di(force_bare), .pad(force_bare_pad) );
    aspida_net_core aspNet ( .nrst(nrst), .clk(clk), .ip_c_req(ip_c_req), 
        .ip_c_we(ip_c_we), .ip_c_mult(ip_c_mult), .ip_c_prd(ip_c_prd), 
        .ip_c_seq(ip_c_seq), .ip_c_ts(ip_c_ts), .ip_c_sel(ip_c_sel), 
        .ip_c_adr(ip_c_adr), .ip_c_dat(ip_c_dat), .ip_c_ack(ip_c_ack), 
        .ip_r_req(ip_r_req), .ip_r_we(ip_r_we), .ip_r_err(ip_r_err), 
        .ip_r_rty(ip_r_rty), .ip_r_acc(ip_r_acc), .ip_r_ts(ip_r_ts), 
        .ip_r_sel(ip_r_sel), .ip_r_dat(ip_r_dat), .ip_r_ack(ip_r_ack), 
        .dp_c_req(dp_c_req), .dp_c_we(dp_c_we), .dp_c_mult(dp_c_mult), 
        .dp_c_prd(dp_c_prd), .dp_c_seq(dp_c_seq), .dp_c_ts(dp_c_ts), 
        .dp_c_sel(dp_c_sel), .dp_c_adr(dp_c_adr), .dp_c_dat(dp_c_dat), 
        .dp_c_ack(dp_c_ack), .dp_r_req(dp_r_req), .dp_r_we(dp_r_we), 
        .dp_r_err(dp_r_err), .dp_r_rty(dp_r_rty), .dp_r_acc(dp_r_acc), 
        .dp_r_ts(dp_r_ts), .dp_r_sel(dp_r_sel), .dp_r_dat(dp_r_dat), 
        .dp_r_ack(dp_r_ack), .ei_c_req(ei_c_req), .ei_c_ack(ei_c_ack), 
        .ei_c_we(ei_c_we), .ei_c_addr({\ei_c_addr[10] , \ei_c_addr[9] , 
        \ei_c_addr[8] , \ei_c_addr[7] , \ei_c_addr[6] , \ei_c_addr[5] , 
        \ei_c_addr[4] , \ei_c_addr[3] , \ei_c_addr[2] , \ei_c_addr[1] , 
        \ei_c_addr[0] }), .ei_r_req(ei_r_req), .ei_r_ack(ei_r_ack), 
        .ei_data_in({\ei_data_in[7] , \ei_data_in[6] , \ei_data_in[5] , 
        \ei_data_in[4] , \ei_data_in[3] , \ei_data_in[2] , \ei_data_in[1] , 
        \ei_data_in[0] }), .ei_data_out({\ei_data_out[7] , \ei_data_out[6] , 
        \ei_data_out[5] , \ei_data_out[4] , \ei_data_out[3] , \ei_data_out[2] , 
        \ei_data_out[1] , \ei_data_out[0] }), .c_BC({\c_BC[4] , \c_BC[3] , 
        \c_BC[2] , \c_BC[1] , \c_BC[0] }), .c_BC_ack(c_BC_ack), .r_BC({
        \r_BC[4] , \r_BC[3] , \r_BC[2] , \r_BC[1] , \r_BC[0] }), .r_BC_ack(
        r_BC_ack), .wish_we_o(wish_we_o), .wish_stb_cyc_o(wish_stb_cyc_o), 
        .wish_ack_i(wish_ack_i), .wish_adr_o({\wish_adr_o[11] , 
        \wish_adr_o[10] , \wish_adr_o[9] , \wish_adr_o[8] , \wish_adr_o[7] , 
        \wish_adr_o[6] , \wish_adr_o[5] , \wish_adr_o[4] , \wish_adr_o[3] , 
        \wish_adr_o[2] , \wish_adr_o[1] , \wish_adr_o[0] }), .wish_dat_i({
        \wish_dat_i[31] , \wish_dat_i[30] , \wish_dat_i[29] , \wish_dat_i[28] , 
        \wish_dat_i[27] , \wish_dat_i[26] , \wish_dat_i[25] , \wish_dat_i[24] , 
        \wish_dat_i[23] , \wish_dat_i[22] , \wish_dat_i[21] , \wish_dat_i[20] , 
        \wish_dat_i[19] , \wish_dat_i[18] , \wish_dat_i[17] , \wish_dat_i[16] , 
        \wish_dat_i[15] , \wish_dat_i[14] , \wish_dat_i[13] , \wish_dat_i[12] , 
        \wish_dat_i[11] , \wish_dat_i[10] , \wish_dat_i[9] , \wish_dat_i[8] , 
        \wish_dat_i[7] , \wish_dat_i[6] , \wish_dat_i[5] , \wish_dat_i[4] , 
        \wish_dat_i[3] , \wish_dat_i[2] , \wish_dat_i[1] , \wish_dat_i[0] }), 
        .wish_dat_o({\wish_dat_o[31] , \wish_dat_o[30] , \wish_dat_o[29] , 
        \wish_dat_o[28] , \wish_dat_o[27] , \wish_dat_o[26] , \wish_dat_o[25] , 
        \wish_dat_o[24] , \wish_dat_o[23] , \wish_dat_o[22] , \wish_dat_o[21] , 
        \wish_dat_o[20] , \wish_dat_o[19] , \wish_dat_o[18] , \wish_dat_o[17] , 
        \wish_dat_o[16] , \wish_dat_o[15] , \wish_dat_o[14] , \wish_dat_o[13] , 
        \wish_dat_o[12] , \wish_dat_o[11] , \wish_dat_o[10] , \wish_dat_o[9] , 
        \wish_dat_o[8] , \wish_dat_o[7] , \wish_dat_o[6] , \wish_dat_o[5] , 
        \wish_dat_o[4] , \wish_dat_o[3] , \wish_dat_o[2] , \wish_dat_o[1] , 
        \wish_dat_o[0] }), .dm_c_req(dm_c_req), .dm_c_we(dm_c_we), .dm_c_mult(
        dm_c_mult), .dm_c_seq(dm_c_seq), .dm_c_prd(dm_c_prd), .dm_c_ts(dm_c_ts
        ), .dm_c_st(dm_c_st), .dm_c_sel(dm_c_sel), .dm_c_adr(dm_c_adr), 
        .dm_c_dat(dm_c_dat), .dm_c_ack(dm_c_ack), .dm_r_req(dm_r_req), 
        .dm_r_err(dm_r_err), .dm_r_rty(dm_r_rty), .dm_r_acc(dm_r_acc), 
        .dm_r_mult(dm_r_mult), .dm_r_ts(dm_r_ts), .dm_r_rt(dm_r_rt), 
        .dm_r_sel(dm_r_sel), .dm_r_dat(dm_r_dat), .dm_r_ack(dm_r_ack), 
        .im_c_req(im_c_req), .im_c_we(im_c_we), .im_c_mult(im_c_mult), 
        .im_c_seq(im_c_seq), .im_c_prd(im_c_prd), .im_c_ts(im_c_ts), .im_c_st(
        im_c_st), .im_c_sel(im_c_sel), .im_c_adr(im_c_adr), .im_c_dat(im_c_dat
        ), .im_c_ack(im_c_ack), .im_r_req(im_r_req), .im_r_err(im_r_err), 
        .im_r_rty(im_r_rty), .im_r_acc(im_r_acc), .im_r_mult(im_r_mult), 
        .im_r_ts(im_r_ts), .im_r_rt(im_r_rt), .im_r_sel(im_r_sel), .im_r_dat(
        im_r_dat), .im_r_ack(im_r_ack), .test_si(test_si), .test_so(test_so), 
        .test_se(test_se), .phi1(phi1), .phi2(phi2), .phi3(phi3), .force_bare(
        force_bare) );
endmodule

