module four_phase_hand(
    input in_ack,
    input in_req,
    input [15:0] in_data,
    input done,

    output out_ack,
    output out_req,
    output [15:0] out_data

);




endmodule