module vmem(clk, addressin,dataout,reset);
input reset;
input clk;
input [14:0] addressin;
output [7:0] dataout;

reg [7:0] dataout;

reg	[7:0]	mem[31:0];
//reg	[7:0]	mem[511:0];

/*reg 	[15:0] i;

initial
begin
	for(i = 0;i< 3072;i = i + 1)
	begin
		mem[i] = i % 8'b11111111;
	end
end*/ 

always @(posedge reset)
begin
// dead //
mem[0]=255;
mem[1]=255;
mem[2]=255;
mem[3]=255;
mem[4]=255;
mem[5]=255;
mem[6]=255;
mem[7]=255;
mem[8]=255;
mem[9]=255;
mem[10]=255;
mem[11]=255;
mem[12]=255;
mem[13]=255;
mem[14]=255;
mem[15]=255;
// live //
mem[16]=0;
mem[17]=0;
mem[18]=0;
mem[19]=0;
mem[20]=0;
mem[21]=0;
mem[22]=0;
mem[23]=0;
mem[24]=0;
mem[25]=0;
mem[26]=0;
mem[27]=0;
mem[28]=0;
mem[29]=0;
mem[30]=0;
mem[31]=0;
/*
mem[0]=255;
mem[1]=255;
mem[2]=255;
mem[3]=255;
mem[4]=255;
mem[5]=255;
mem[6]=255;
mem[7]=255;
mem[8]=255;
mem[9]=255;
mem[10]=255;
mem[11]=255;
mem[12]=255;
mem[13]=255;
mem[14]=255;
mem[15]=255;
mem[16]=0;
mem[17]=0;
mem[18]=0;
mem[19]=0;
mem[20]=0;
mem[21]=0;
mem[22]=0;
mem[23]=0;
mem[24]=0;
mem[25]=0;
mem[26]=0;
mem[27]=0;
mem[28]=0;
mem[29]=0;
mem[30]=0;
mem[31]=0;
mem[32]=1;
mem[33]=1;
mem[34]=1;
mem[35]=1;
mem[36]=1;
mem[37]=1;
mem[38]=1;
mem[39]=0;
mem[40]=1;
mem[41]=1;
mem[42]=1;
mem[43]=1;
mem[44]=1;
mem[45]=1;
mem[46]=1;
mem[47]=1;
mem[48]=1;
mem[49]=1;
mem[50]=1;
mem[51]=1;
mem[52]=1;
mem[53]=1;
mem[54]=1;
mem[55]=1;
mem[56]=1;
mem[57]=1;
mem[58]=1;
mem[59]=0;
mem[60]=1;
mem[61]=1;
mem[62]=1;
mem[63]=1;
mem[64]=1;
mem[65]=1;
mem[66]=1;
mem[67]=1;
mem[68]=1;
mem[69]=1;
mem[70]=1;
mem[71]=1;
mem[72]=1;
mem[73]=1;
mem[74]=1;
mem[75]=1;
mem[76]=1;
mem[77]=1;
mem[78]=1;
mem[79]=1;
mem[80]=1;
mem[81]=1;
mem[82]=1;
mem[83]=1;
mem[84]=1;
mem[85]=1;
mem[86]=1;
mem[87]=1;
mem[88]=1;
mem[89]=1;
mem[90]=1;
mem[91]=1;
mem[92]=1;
mem[93]=1;
mem[94]=1;
mem[95]=1;
mem[96]=1;
mem[97]=1;
mem[98]=1;
mem[99]=1;
mem[100]=1;
mem[101]=1;
mem[102]=1;
mem[103]=1;
mem[104]=1;
mem[105]=1;
mem[106]=1;
mem[107]=1;
mem[108]=1;
mem[109]=1;
mem[110]=1;
mem[111]=1;
mem[112]=1;
mem[113]=1;
mem[114]=1;
mem[115]=1;
mem[116]=1;
mem[117]=1;
mem[118]=1;
mem[119]=1;
mem[120]=1;
mem[121]=1;
mem[122]=1;
mem[123]=1;
mem[124]=1;
mem[125]=1;
mem[126]=1;
mem[127]=1;
mem[128]=1;
mem[129]=0;
mem[130]=0;
mem[131]=0;
mem[132]=0;
mem[133]=255;
mem[134]=255;
mem[135]=0;
mem[136]=0;
mem[137]=255;
mem[138]=255;
mem[139]=0;
mem[140]=0;
mem[141]=0;
mem[142]=0;
mem[143]=0;
mem[144]=0;
mem[145]=250;
mem[146]=250;
mem[147]=250;
mem[148]=250;
mem[149]=250;
mem[150]=0;
mem[151]=0;
mem[152]=250;
mem[153]=250;
mem[154]=0;
mem[155]=0;
mem[156]=250;
mem[157]=250;
mem[158]=250;
mem[159]=250;
mem[160]=250;
mem[161]=1;
mem[162]=0;
mem[163]=1;
mem[164]=0;
mem[165]=1;
mem[166]=0;
mem[167]=1;
mem[168]=0;
mem[169]=1;
mem[170]=0;
mem[171]=1;
mem[172]=0;
mem[173]=1;
mem[174]=0;
mem[175]=1;
mem[176]=0;
mem[177]=1;
mem[178]=0;
mem[179]=1;
mem[180]=0;
mem[181]=1;
mem[182]=0;
mem[183]=1;
mem[184]=0;
mem[185]=1;
mem[186]=0;
mem[187]=1;
mem[188]=0;
mem[189]=1;
mem[190]=150;
mem[191]=1;
mem[192]=0;
mem[193]=1;
mem[194]=0;
mem[195]=1;
mem[196]=0;
mem[197]=1;
mem[198]=0;
mem[199]=1;
mem[200]=0;
mem[201]=1;
mem[202]=0;
mem[203]=1;
mem[204]=0;
mem[205]=1;
mem[206]=0;
mem[207]=1;
mem[208]=0;
mem[209]=1;
mem[210]=0;
mem[211]=1;
mem[212]=0;
mem[213]=1;
mem[214]=0;
mem[215]=1;
mem[216]=0;
mem[217]=1;
mem[218]=0;
mem[219]=1;
mem[220]=0;
mem[221]=1;
mem[222]=0;
mem[223]=1;
mem[224]=0;
mem[225]=1;
mem[226]=0;
mem[227]=1;
mem[228]=0;
mem[229]=1;
mem[230]=0;
mem[231]=1;
mem[232]=0;
mem[233]=1;
mem[234]=0;
mem[235]=1;
mem[236]=0;
mem[237]=1;
mem[238]=0;
mem[239]=1;
mem[240]=0;
mem[241]=1;
mem[242]=0;
mem[243]=1;
mem[244]=0;
mem[245]=1;
mem[246]=0;
mem[247]=1;
mem[248]=0;
mem[249]=1;
mem[250]=0;
mem[251]=1;
mem[252]=0;
mem[253]=1;
mem[254]=0;
mem[255]=1;
mem[256]=0;
mem[257]=0;
mem[258]=0;
mem[259]=0;
mem[260]=0;
mem[261]=0;
mem[262]=0;
mem[263]=0;
mem[264]=0;
mem[265]=0;
mem[266]=0;
mem[267]=0;
mem[268]=0;
mem[269]=0;
mem[270]=0;
mem[271]=0;
mem[272]=0;
mem[273]=0;
mem[274]=0;
mem[275]=0;
mem[276]=0;
mem[277]=0;
mem[278]=0;
mem[279]=0;
mem[280]=0;
mem[281]=0;
mem[282]=0;
mem[283]=0;
mem[284]=0;
mem[285]=0;
mem[286]=0;
mem[287]=0;
mem[288]=0;
mem[289]=0;
mem[290]=0;
mem[291]=0;
mem[292]=0;
mem[293]=0;
mem[294]=0;
mem[295]=0;
mem[296]=0;
mem[297]=0;
mem[298]=0;
mem[299]=0;
mem[300]=0;
mem[301]=0;
mem[302]=0;
mem[303]=0;
mem[304]=0;
mem[305]=0;
mem[306]=0;
mem[307]=0;
mem[308]=0;
mem[309]=0;
mem[310]=0;
mem[311]=0;
mem[312]=0;
mem[313]=0;
mem[314]=0;
mem[315]=0;
mem[316]=0;
mem[317]=0;
mem[318]=0;
mem[319]=0;
mem[320]=0;
mem[321]=0;
mem[322]=0;
mem[323]=0;
mem[324]=0;
mem[325]=0;
mem[326]=0;
mem[327]=0;
mem[328]=0;
mem[329]=0;
mem[330]=0;
mem[331]=0;
mem[332]=0;
mem[333]=0;
mem[334]=0;
mem[335]=0;
mem[336]=0;
mem[337]=0;
mem[338]=0;
mem[339]=0;
mem[340]=0;
mem[341]=0;
mem[342]=0;
mem[343]=0;
mem[344]=0;
mem[345]=0;
mem[346]=0;
mem[347]=0;
mem[348]=0;
mem[349]=0;
mem[350]=0;
mem[351]=0;
mem[352]=0;
mem[353]=0;
mem[354]=0;
mem[355]=0;
mem[356]=0;
mem[357]=0;
mem[358]=0;
mem[359]=0;
mem[360]=0;
mem[361]=0;
mem[362]=0;
mem[363]=0;
mem[364]=0;
mem[365]=0;
mem[366]=0;
mem[367]=0;
mem[368]=0;
mem[369]=0;
mem[370]=0;
mem[371]=0;
mem[372]=0;
mem[373]=0;
mem[374]=0;
mem[375]=0;
mem[376]=0;
mem[377]=0;
mem[378]=0;
mem[379]=0;
mem[380]=0;
mem[381]=0;
mem[382]=0;
mem[383]=0;
mem[384]=0;
mem[385]=0;
mem[386]=0;
mem[387]=0;
mem[388]=0;
mem[389]=0;
mem[390]=0;
mem[391]=0;
mem[392]=0;
mem[393]=0;
mem[394]=0;
mem[395]=0;
mem[396]=0;
mem[397]=0;
mem[398]=0;
mem[399]=0;
mem[400]=0;
mem[401]=0;
mem[402]=0;
mem[403]=0;
mem[404]=0;
mem[405]=0;
mem[406]=0;
mem[407]=0;
mem[408]=0;
mem[409]=0;
mem[410]=0;
mem[411]=0;
mem[412]=0;
mem[413]=0;
mem[414]=0;
mem[415]=0;
mem[416]=0;
mem[417]=0;
mem[418]=0;
mem[419]=0;
mem[420]=0;
mem[421]=0;
mem[422]=0;
mem[423]=0;
mem[424]=0;
mem[425]=0;
mem[426]=0;
mem[427]=0;
mem[428]=0;
mem[429]=0;
mem[430]=0;
mem[431]=0;
mem[432]=0;
mem[433]=0;
mem[434]=0;
mem[435]=0;
mem[436]=0;
mem[437]=0;
mem[438]=0;
mem[439]=0;
mem[440]=0;
mem[441]=0;
mem[442]=0;
mem[443]=0;
mem[444]=0;
mem[445]=0;
mem[446]=0;
mem[447]=0;
mem[448]=0;
mem[449]=0;
mem[450]=0;
mem[451]=0;
mem[452]=0;
mem[453]=0;
mem[454]=0;
mem[455]=0;
mem[456]=0;
mem[457]=0;
mem[458]=0;
mem[459]=0;
mem[460]=0;
mem[461]=0;
mem[462]=0;
mem[463]=0;
mem[464]=0;
mem[465]=0;
mem[466]=0;
mem[467]=0;
mem[468]=0;
mem[469]=0;
mem[470]=0;
mem[471]=0;
mem[472]=0;
mem[473]=0;
mem[474]=0;
mem[475]=0;
mem[476]=0;
mem[477]=0;
mem[478]=0;
mem[479]=0;
mem[480]=0;
mem[481]=0;
mem[482]=0;
mem[483]=0;
mem[484]=0;
mem[485]=0;
mem[486]=0;
mem[487]=0;
mem[488]=0;
mem[489]=0;
mem[490]=0;
mem[491]=0;
mem[492]=0;
mem[493]=0;
mem[494]=0;
mem[495]=0;
mem[496]=0;
mem[497]=0;
mem[498]=0;
mem[499]=0;
mem[500]=0;
mem[501]=0;
mem[502]=0;
mem[503]=0;
mem[504]=0;
mem[505]=0;
mem[506]=0;
mem[507]=0;
mem[508]=0;
mem[509]=0;
mem[510]=0;
mem[511]=0;
*/
end	

//always @(addressin)
always @(posedge clk)
begin
	dataout = mem[addressin];
end

endmodule
